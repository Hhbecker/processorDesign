<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-13.7483,62.4001,490.92,-218.252</PageViewport>
<gate>
<ID>389</ID>
<type>DA_FROM</type>
<position>385.5,-99</position>
<input>
<ID>IN_0</ID>531 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load bit 4 (DR)</lparam></gate>
<gate>
<ID>391</ID>
<type>AA_MUX_2x1</type>
<position>138,-143</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>480 </output>
<input>
<ID>SEL_0</ID>462 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_MUX_2x1</type>
<position>205.5,-128</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>460 </input>
<output>
<ID>OUT</ID>463 </output>
<input>
<ID>SEL_0</ID>462 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>395</ID>
<type>DE_TO</type>
<position>225.5,56</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load bit 4 (DR)</lparam></gate>
<gate>
<ID>396</ID>
<type>AA_MUX_2x1</type>
<position>111,-149</position>
<input>
<ID>IN_0</ID>479 </input>
<input>
<ID>IN_1</ID>476 </input>
<output>
<ID>OUT</ID>482 </output>
<input>
<ID>SEL_0</ID>462 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>397</ID>
<type>AA_MUX_2x1</type>
<position>165,-137</position>
<input>
<ID>IN_0</ID>470 </input>
<input>
<ID>IN_1</ID>466 </input>
<output>
<ID>OUT</ID>469 </output>
<input>
<ID>SEL_0</ID>462 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>398</ID>
<type>AA_TOGGLE</type>
<position>290.5,42.5</position>
<output>
<ID>OUT_0</ID>739 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>402</ID>
<type>AA_MUX_2x1</type>
<position>124.5,-146</position>
<input>
<ID>IN_0</ID>478 </input>
<input>
<ID>IN_1</ID>475 </input>
<output>
<ID>OUT</ID>481 </output>
<input>
<ID>SEL_0</ID>462 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>403</ID>
<type>AA_MUX_2x1</type>
<position>191.5,-131</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>459 </input>
<output>
<ID>OUT</ID>465 </output>
<input>
<ID>SEL_0</ID>462 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>404</ID>
<type>DA_FROM</type>
<position>139.5,-108</position>
<input>
<ID>IN_0</ID>430 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt5</lparam></gate>
<gate>
<ID>406</ID>
<type>DA_FROM</type>
<position>190.5,-108</position>
<input>
<ID>IN_0</ID>451 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt2</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_TOGGLE</type>
<position>293.5,42.5</position>
<output>
<ID>OUT_0</ID>740 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>410</ID>
<type>DA_FROM</type>
<position>142.5,-108</position>
<input>
<ID>IN_0</ID>429 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt4</lparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>107,-124</position>
<input>
<ID>IN_0</ID>479 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp7</lparam></gate>
<gate>
<ID>413</ID>
<type>DA_FROM</type>
<position>134,-126</position>
<input>
<ID>IN_0</ID>477 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp5</lparam></gate>
<gate>
<ID>414</ID>
<type>DA_FROM</type>
<position>147.5,-125</position>
<input>
<ID>IN_0</ID>471 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp4</lparam></gate>
<gate>
<ID>416</ID>
<type>DA_FROM</type>
<position>286,51</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Load</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>184.5,-108</position>
<input>
<ID>IN_0</ID>454 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut0</lparam></gate>
<gate>
<ID>418</ID>
<type>DA_FROM</type>
<position>193.5,-108</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt1</lparam></gate>
<gate>
<ID>420</ID>
<type>DA_FROM</type>
<position>289,48</position>
<input>
<ID>IN_0</ID>739 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID CEnable</lparam></gate>
<gate>
<ID>422</ID>
<type>DA_FROM</type>
<position>201.5,-125</position>
<input>
<ID>IN_0</ID>461 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID PCUp0</lparam></gate>
<gate>
<ID>423</ID>
<type>DA_FROM</type>
<position>187.5,-108</position>
<input>
<ID>IN_0</ID>450 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt3</lparam></gate>
<gate>
<ID>425</ID>
<type>DA_FROM</type>
<position>136.5,-108</position>
<input>
<ID>IN_0</ID>431 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt6</lparam></gate>
<gate>
<ID>426</ID>
<type>AA_TOGGLE</type>
<position>297.5,25.5</position>
<output>
<ID>OUT_0</ID>741 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>427</ID>
<type>DA_FROM</type>
<position>196.5,-108</position>
<input>
<ID>IN_0</ID>453 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt0</lparam></gate>
<gate>
<ID>428</ID>
<type>DA_FROM</type>
<position>188,-126</position>
<input>
<ID>IN_0</ID>464 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID PCUp1</lparam></gate>
<gate>
<ID>429</ID>
<type>DA_FROM</type>
<position>174.5,-125</position>
<input>
<ID>IN_0</ID>467 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID PCUp2</lparam></gate>
<gate>
<ID>430</ID>
<type>DA_FROM</type>
<position>120.5,-125</position>
<input>
<ID>IN_0</ID>478 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp6</lparam></gate>
<gate>
<ID>431</ID>
<type>DA_FROM</type>
<position>161,-124</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp3</lparam></gate>
<gate>
<ID>432</ID>
<type>DE_TO</type>
<position>178.5,-154</position>
<input>
<ID>IN_0</ID>468 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux2</lparam></gate>
<gate>
<ID>433</ID>
<type>DE_TO</type>
<position>165,-154</position>
<input>
<ID>IN_0</ID>469 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux3</lparam></gate>
<gate>
<ID>434</ID>
<type>DE_TO</type>
<position>151.5,-154</position>
<input>
<ID>IN_0</ID>473 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux4</lparam></gate>
<gate>
<ID>435</ID>
<type>DE_TO</type>
<position>111,-154</position>
<input>
<ID>IN_0</ID>482 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux7</lparam></gate>
<gate>
<ID>436</ID>
<type>DE_TO</type>
<position>205.5,-154</position>
<input>
<ID>IN_0</ID>463 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux0</lparam></gate>
<gate>
<ID>437</ID>
<type>DE_TO</type>
<position>191.5,-154</position>
<input>
<ID>IN_0</ID>465 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux1</lparam></gate>
<gate>
<ID>438</ID>
<type>DE_TO</type>
<position>124.5,-154</position>
<input>
<ID>IN_0</ID>481 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux6</lparam></gate>
<gate>
<ID>439</ID>
<type>DE_TO</type>
<position>138,-154</position>
<input>
<ID>IN_0</ID>480 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux5</lparam></gate>
<gate>
<ID>440</ID>
<type>DA_FROM</type>
<position>133.5,-108</position>
<input>
<ID>IN_0</ID>448 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt7</lparam></gate>
<gate>
<ID>441</ID>
<type>DA_FROM</type>
<position>178.5,-108</position>
<input>
<ID>IN_0</ID>456 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut2</lparam></gate>
<gate>
<ID>442</ID>
<type>DA_FROM</type>
<position>130.5,-108</position>
<input>
<ID>IN_0</ID>425 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut4</lparam></gate>
<gate>
<ID>443</ID>
<type>DA_FROM</type>
<position>124.5,-108</position>
<input>
<ID>IN_0</ID>427 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut6</lparam></gate>
<gate>
<ID>444</ID>
<type>DA_FROM</type>
<position>175.5,-108</position>
<input>
<ID>IN_0</ID>457 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut3</lparam></gate>
<gate>
<ID>445</ID>
<type>DA_FROM</type>
<position>127.5,-108</position>
<input>
<ID>IN_0</ID>426 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut5</lparam></gate>
<gate>
<ID>446</ID>
<type>DA_FROM</type>
<position>121.5,-108</position>
<input>
<ID>IN_0</ID>428 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut7</lparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>181.5,-108</position>
<input>
<ID>IN_0</ID>455 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut1</lparam></gate>
<gate>
<ID>448</ID>
<type>DA_FROM</type>
<position>365.5,-55.5</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>449</ID>
<type>AA_TOGGLE</type>
<position>240,11.5</position>
<output>
<ID>OUT_0</ID>742 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>450</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>377,-36.5</position>
<input>
<ID>ENABLE_0</ID>683 </input>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>485 </input>
<input>
<ID>IN_2</ID>486 </input>
<input>
<ID>IN_3</ID>487 </input>
<input>
<ID>IN_4</ID>488 </input>
<input>
<ID>IN_5</ID>489 </input>
<input>
<ID>IN_6</ID>490 </input>
<input>
<ID>IN_7</ID>491 </input>
<output>
<ID>OUT_0</ID>631 </output>
<output>
<ID>OUT_1</ID>630 </output>
<output>
<ID>OUT_2</ID>629 </output>
<output>
<ID>OUT_3</ID>628 </output>
<output>
<ID>OUT_4</ID>627 </output>
<output>
<ID>OUT_5</ID>626 </output>
<output>
<ID>OUT_6</ID>597 </output>
<output>
<ID>OUT_7</ID>640 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>451</ID>
<type>DA_FROM</type>
<position>366,-47.5</position>
<input>
<ID>IN_0</ID>485 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>452</ID>
<type>DA_FROM</type>
<position>363.5,-42.5</position>
<input>
<ID>IN_0</ID>486 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>453</ID>
<type>AA_LABEL</type>
<position>519.5,61.5</position>
<gparam>LABEL_TEXT Register File</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>454</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>657,-62</position>
<input>
<ID>IN_0</ID>730 </input>
<input>
<ID>IN_1</ID>736 </input>
<input>
<ID>IN_2</ID>507 </input>
<input>
<ID>IN_3</ID>505 </input>
<input>
<ID>IN_4</ID>503 </input>
<input>
<ID>IN_5</ID>501 </input>
<input>
<ID>IN_6</ID>668 </input>
<input>
<ID>IN_7</ID>641 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>455</ID>
<type>DE_TO</type>
<position>670.5,-17.5</position>
<input>
<ID>IN_0</ID>596 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>456</ID>
<type>DE_TO</type>
<position>670,-24.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>457</ID>
<type>DE_TO</type>
<position>670,-27.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>458</ID>
<type>DE_TO</type>
<position>670,-31</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>459</ID>
<type>DE_TO</type>
<position>670.5,-34</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>460</ID>
<type>DE_TO</type>
<position>670.5,-37</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>461</ID>
<type>DE_TO</type>
<position>671,-40.5</position>
<input>
<ID>IN_0</ID>729 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>462</ID>
<type>DE_TO</type>
<position>670,-21.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>463</ID>
<type>DE_TO</type>
<position>672.5,-55.5</position>
<input>
<ID>IN_0</ID>641 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>464</ID>
<type>DA_FROM</type>
<position>361.5,-37</position>
<input>
<ID>IN_0</ID>487 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>465</ID>
<type>DA_FROM</type>
<position>344.5,-33</position>
<input>
<ID>IN_0</ID>488 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>466</ID>
<type>DA_FROM</type>
<position>345.5,-27.5</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>467</ID>
<type>DA_FROM</type>
<position>345,-23.5</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>468</ID>
<type>DA_FROM</type>
<position>345,-19.5</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>469</ID>
<type>DE_TO</type>
<position>673,-79</position>
<input>
<ID>IN_0</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>470</ID>
<type>AE_REGISTER8</type>
<position>144,-31</position>
<input>
<ID>IN_0</ID>584 </input>
<input>
<ID>IN_1</ID>585 </input>
<input>
<ID>IN_2</ID>586 </input>
<input>
<ID>IN_3</ID>587 </input>
<input>
<ID>IN_4</ID>588 </input>
<input>
<ID>IN_5</ID>589 </input>
<input>
<ID>IN_6</ID>590 </input>
<input>
<ID>IN_7</ID>591 </input>
<output>
<ID>OUT_0</ID>534 </output>
<output>
<ID>OUT_1</ID>533 </output>
<output>
<ID>OUT_2</ID>499 </output>
<output>
<ID>OUT_3</ID>498 </output>
<output>
<ID>OUT_4</ID>497 </output>
<output>
<ID>OUT_5</ID>496 </output>
<output>
<ID>OUT_6</ID>495 </output>
<output>
<ID>OUT_7</ID>494 </output>
<input>
<ID>clear</ID>492 </input>
<input>
<ID>clock</ID>642 </input>
<input>
<ID>load</ID>535 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>471</ID>
<type>DE_TO</type>
<position>672.5,-58.5</position>
<input>
<ID>IN_0</ID>668 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>472</ID>
<type>AA_LABEL</type>
<position>302,85.5</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>473</ID>
<type>AA_LABEL</type>
<position>151.5,-90</position>
<gparam>LABEL_TEXT PC adder for offset in Branch Case</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>474</ID>
<type>DE_TO</type>
<position>672.5,-62.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>475</ID>
<type>DE_TO</type>
<position>672.5,-66.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>476</ID>
<type>DE_TO</type>
<position>673.5,-75.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>477</ID>
<type>DE_TO</type>
<position>673,-70.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>478</ID>
<type>DE_TO</type>
<position>673.5,-73</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>479</ID>
<type>AE_REGISTER8</type>
<position>198.5,55</position>
<input>
<ID>IN_0</ID>639 </input>
<input>
<ID>IN_1</ID>638 </input>
<input>
<ID>IN_2</ID>637 </input>
<input>
<ID>IN_3</ID>636 </input>
<input>
<ID>IN_4</ID>635 </input>
<input>
<ID>IN_5</ID>634 </input>
<input>
<ID>IN_6</ID>633 </input>
<input>
<ID>IN_7</ID>632 </input>
<output>
<ID>OUT_0</ID>545 </output>
<output>
<ID>OUT_1</ID>544 </output>
<output>
<ID>OUT_2</ID>543 </output>
<output>
<ID>OUT_3</ID>542 </output>
<output>
<ID>OUT_4</ID>541 </output>
<output>
<ID>OUT_5</ID>540 </output>
<output>
<ID>OUT_6</ID>539 </output>
<output>
<ID>OUT_7</ID>538 </output>
<input>
<ID>clear</ID>546 </input>
<input>
<ID>clock</ID>642 </input>
<input>
<ID>load</ID>547 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>480</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>205.5,55.5</position>
<input>
<ID>ENABLE_0</ID>673 </input>
<input>
<ID>IN_0</ID>545 </input>
<input>
<ID>IN_1</ID>544 </input>
<input>
<ID>IN_2</ID>543 </input>
<input>
<ID>IN_3</ID>542 </input>
<input>
<ID>IN_4</ID>541 </input>
<input>
<ID>IN_5</ID>540 </input>
<input>
<ID>IN_6</ID>539 </input>
<input>
<ID>IN_7</ID>538 </input>
<output>
<ID>OUT_0</ID>675 </output>
<output>
<ID>OUT_1</ID>676 </output>
<output>
<ID>OUT_2</ID>677 </output>
<output>
<ID>OUT_3</ID>678 </output>
<output>
<ID>OUT_4</ID>738 </output>
<output>
<ID>OUT_5</ID>660 </output>
<output>
<ID>OUT_6</ID>671 </output>
<output>
<ID>OUT_7</ID>672 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>481</ID>
<type>AA_TOGGLE</type>
<position>199.5,44</position>
<output>
<ID>OUT_0</ID>546 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>482</ID>
<type>AA_TOGGLE</type>
<position>415,30.5</position>
<output>
<ID>OUT_0</ID>595 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>483</ID>
<type>AA_LABEL</type>
<position>205,44.5</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>484</ID>
<type>AA_LABEL</type>
<position>197,71</position>
<gparam>LABEL_TEXT Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>485</ID>
<type>AA_TOGGLE</type>
<position>415,35</position>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>486</ID>
<type>AA_LABEL</type>
<position>211,71</position>
<gparam>LABEL_TEXT IR control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>487</ID>
<type>AA_LABEL</type>
<position>207,76.5</position>
<gparam>LABEL_TEXT Instruction Register</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>488</ID>
<type>AA_TOGGLE</type>
<position>143,-39.5</position>
<output>
<ID>OUT_0</ID>492 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>489</ID>
<type>AA_LABEL</type>
<position>143.5,-42</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>490</ID>
<type>AA_LABEL</type>
<position>656,-14</position>
<gparam>LABEL_TEXT SR1 Out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>491</ID>
<type>AA_TOGGLE</type>
<position>413.5,45.5</position>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>492</ID>
<type>AA_LABEL</type>
<position>657,-51</position>
<gparam>LABEL_TEXT SR2 Out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>493</ID>
<type>AA_LABEL</type>
<position>118,2</position>
<gparam>LABEL_TEXT Memory</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>494</ID>
<type>AE_RAM_8x8</type>
<position>126.5,-18</position>
<input>
<ID>ADDRESS_0</ID>555 </input>
<input>
<ID>ADDRESS_1</ID>554 </input>
<input>
<ID>ADDRESS_2</ID>553 </input>
<input>
<ID>ADDRESS_3</ID>552 </input>
<input>
<ID>ADDRESS_4</ID>551 </input>
<input>
<ID>ADDRESS_5</ID>550 </input>
<input>
<ID>ADDRESS_6</ID>549 </input>
<input>
<ID>ADDRESS_7</ID>548 </input>
<input>
<ID>DATA_IN_0</ID>584 </input>
<input>
<ID>DATA_IN_1</ID>585 </input>
<input>
<ID>DATA_IN_2</ID>586 </input>
<input>
<ID>DATA_IN_3</ID>587 </input>
<input>
<ID>DATA_IN_4</ID>588 </input>
<input>
<ID>DATA_IN_5</ID>589 </input>
<input>
<ID>DATA_IN_6</ID>590 </input>
<input>
<ID>DATA_IN_7</ID>591 </input>
<output>
<ID>DATA_OUT_0</ID>584 </output>
<output>
<ID>DATA_OUT_1</ID>585 </output>
<output>
<ID>DATA_OUT_2</ID>586 </output>
<output>
<ID>DATA_OUT_3</ID>587 </output>
<output>
<ID>DATA_OUT_4</ID>588 </output>
<output>
<ID>DATA_OUT_5</ID>589 </output>
<output>
<ID>DATA_OUT_6</ID>590 </output>
<output>
<ID>DATA_OUT_7</ID>591 </output>
<input>
<ID>ENABLE_0</ID>743 </input>
<input>
<ID>write_clock</ID>642 </input>
<input>
<ID>write_enable</ID>592 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>495</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>157.5,-30.5</position>
<input>
<ID>ENABLE_0</ID>493 </input>
<input>
<ID>IN_0</ID>534 </input>
<input>
<ID>IN_1</ID>533 </input>
<input>
<ID>IN_2</ID>499 </input>
<input>
<ID>IN_3</ID>498 </input>
<input>
<ID>IN_4</ID>497 </input>
<input>
<ID>IN_5</ID>496 </input>
<input>
<ID>IN_6</ID>495 </input>
<input>
<ID>IN_7</ID>494 </input>
<output>
<ID>OUT_0</ID>607 </output>
<output>
<ID>OUT_1</ID>606 </output>
<output>
<ID>OUT_2</ID>605 </output>
<output>
<ID>OUT_3</ID>604 </output>
<output>
<ID>OUT_4</ID>603 </output>
<output>
<ID>OUT_5</ID>602 </output>
<output>
<ID>OUT_6</ID>601 </output>
<output>
<ID>OUT_7</ID>600 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>496</ID>
<type>DA_FROM</type>
<position>143.5,-22.5</position>
<input>
<ID>IN_0</ID>535 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRload</lparam></gate>
<gate>
<ID>497</ID>
<type>DA_FROM</type>
<position>160.5,-23</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID MDRsend</lparam></gate>
<gate>
<ID>498</ID>
<type>AE_REGISTER8</type>
<position>290.5,32.5</position>
<input>
<ID>IN_0</ID>563 </input>
<input>
<ID>IN_1</ID>562 </input>
<input>
<ID>IN_2</ID>561 </input>
<input>
<ID>IN_3</ID>560 </input>
<input>
<ID>IN_4</ID>559 </input>
<input>
<ID>IN_5</ID>558 </input>
<input>
<ID>IN_6</ID>557 </input>
<input>
<ID>IN_7</ID>556 </input>
<output>
<ID>OUT_0</ID>570 </output>
<output>
<ID>OUT_1</ID>571 </output>
<output>
<ID>OUT_2</ID>572 </output>
<output>
<ID>OUT_3</ID>569 </output>
<output>
<ID>OUT_4</ID>565 </output>
<output>
<ID>OUT_5</ID>566 </output>
<output>
<ID>OUT_6</ID>567 </output>
<output>
<ID>OUT_7</ID>568 </output>
<input>
<ID>clear</ID>741 </input>
<input>
<ID>clock</ID>642 </input>
<input>
<ID>count_enable</ID>739 </input>
<input>
<ID>count_up</ID>740 </input>
<input>
<ID>load</ID>564 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>499</ID>
<type>AA_LABEL</type>
<position>278,61.5</position>
<gparam>LABEL_TEXT CountIn</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>500</ID>
<type>AA_TOGGLE</type>
<position>282.5,61</position>
<output>
<ID>OUT_0</ID>574 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>501</ID>
<type>AA_TOGGLE</type>
<position>287.5,42.5</position>
<output>
<ID>OUT_0</ID>564 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>502</ID>
<type>DA_FROM</type>
<position>279.5,43.5</position>
<input>
<ID>IN_0</ID>556 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux7</lparam></gate>
<gate>
<ID>503</ID>
<type>DA_FROM</type>
<position>279.5,40.5</position>
<input>
<ID>IN_0</ID>557 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux6</lparam></gate>
<gate>
<ID>504</ID>
<type>DA_FROM</type>
<position>279.5,37.5</position>
<input>
<ID>IN_0</ID>558 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux5</lparam></gate>
<gate>
<ID>505</ID>
<type>DA_FROM</type>
<position>279.5,34.5</position>
<input>
<ID>IN_0</ID>559 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux4</lparam></gate>
<gate>
<ID>506</ID>
<type>DA_FROM</type>
<position>279.5,31.5</position>
<input>
<ID>IN_0</ID>560 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux3</lparam></gate>
<gate>
<ID>507</ID>
<type>DA_FROM</type>
<position>279.5,28.5</position>
<input>
<ID>IN_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux2</lparam></gate>
<gate>
<ID>508</ID>
<type>DA_FROM</type>
<position>279.5,25.5</position>
<input>
<ID>IN_0</ID>562 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux1</lparam></gate>
<gate>
<ID>509</ID>
<type>DA_FROM</type>
<position>279.5,22.5</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux0</lparam></gate>
<gate>
<ID>510</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>318.5,33</position>
<input>
<ID>ENABLE_0</ID>651 </input>
<input>
<ID>IN_0</ID>570 </input>
<input>
<ID>IN_1</ID>571 </input>
<input>
<ID>IN_2</ID>572 </input>
<input>
<ID>IN_3</ID>569 </input>
<input>
<ID>IN_4</ID>565 </input>
<input>
<ID>IN_5</ID>566 </input>
<input>
<ID>IN_6</ID>567 </input>
<input>
<ID>IN_7</ID>568 </input>
<output>
<ID>OUT_0</ID>649 </output>
<output>
<ID>OUT_1</ID>650 </output>
<output>
<ID>OUT_2</ID>652 </output>
<output>
<ID>OUT_3</ID>653 </output>
<output>
<ID>OUT_4</ID>654 </output>
<output>
<ID>OUT_5</ID>655 </output>
<output>
<ID>OUT_6</ID>656 </output>
<output>
<ID>OUT_7</ID>657 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>511</ID>
<type>DE_TO</type>
<position>309,71</position>
<input>
<ID>IN_0</ID>580 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp1</lparam></gate>
<gate>
<ID>512</ID>
<type>DE_TO</type>
<position>312,71</position>
<input>
<ID>IN_0</ID>581 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp2</lparam></gate>
<gate>
<ID>513</ID>
<type>DE_TO</type>
<position>315,71</position>
<input>
<ID>IN_0</ID>582 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp3</lparam></gate>
<gate>
<ID>514</ID>
<type>DE_TO</type>
<position>289,71</position>
<input>
<ID>IN_0</ID>576 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp4</lparam></gate>
<gate>
<ID>515</ID>
<type>DE_TO</type>
<position>306,71</position>
<input>
<ID>IN_0</ID>583 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp0</lparam></gate>
<gate>
<ID>516</ID>
<type>DE_TO</type>
<position>292,71</position>
<input>
<ID>IN_0</ID>577 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp5</lparam></gate>
<gate>
<ID>517</ID>
<type>DE_TO</type>
<position>298,71</position>
<input>
<ID>IN_0</ID>579 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp7</lparam></gate>
<gate>
<ID>518</ID>
<type>DE_TO</type>
<position>295,71</position>
<input>
<ID>IN_0</ID>578 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp6</lparam></gate>
<gate>
<ID>519</ID>
<type>AA_TOGGLE</type>
<position>414,49</position>
<output>
<ID>OUT_0</ID>528 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>520</ID>
<type>AE_FULLADDER_4BIT</type>
<position>293.5,62</position>
<input>
<ID>IN_0</ID>565 </input>
<input>
<ID>IN_1</ID>566 </input>
<input>
<ID>IN_2</ID>567 </input>
<input>
<ID>IN_3</ID>568 </input>
<output>
<ID>OUT_0</ID>576 </output>
<output>
<ID>OUT_1</ID>577 </output>
<output>
<ID>OUT_2</ID>578 </output>
<output>
<ID>OUT_3</ID>579 </output>
<input>
<ID>carry_in</ID>574 </input>
<output>
<ID>carry_out</ID>573 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>521</ID>
<type>AE_FULLADDER_4BIT</type>
<position>310.5,62</position>
<input>
<ID>IN_0</ID>570 </input>
<input>
<ID>IN_1</ID>571 </input>
<input>
<ID>IN_2</ID>572 </input>
<input>
<ID>IN_3</ID>569 </input>
<output>
<ID>OUT_0</ID>583 </output>
<output>
<ID>OUT_1</ID>580 </output>
<output>
<ID>OUT_2</ID>581 </output>
<output>
<ID>OUT_3</ID>582 </output>
<input>
<ID>carry_in</ID>573 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>522</ID>
<type>AA_LABEL</type>
<position>305.5,39</position>
<gparam>LABEL_TEXT PCOut</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>523</ID>
<type>DE_TO</type>
<position>230.5,-35.5</position>
<input>
<ID>IN_0</ID>536 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRsend</lparam></gate>
<gate>
<ID>524</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>119.5,-44</position>
<input>
<ID>ENABLE_0</ID>592 </input>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>598 </input>
<input>
<ID>IN_2</ID>647 </input>
<input>
<ID>IN_3</ID>648 </input>
<input>
<ID>IN_4</ID>645 </input>
<input>
<ID>IN_5</ID>644 </input>
<input>
<ID>IN_6</ID>643 </input>
<input>
<ID>IN_7</ID>593 </input>
<output>
<ID>OUT_0</ID>584 </output>
<output>
<ID>OUT_1</ID>585 </output>
<output>
<ID>OUT_2</ID>586 </output>
<output>
<ID>OUT_3</ID>587 </output>
<output>
<ID>OUT_4</ID>588 </output>
<output>
<ID>OUT_5</ID>589 </output>
<output>
<ID>OUT_6</ID>590 </output>
<output>
<ID>OUT_7</ID>591 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>525</ID>
<type>AA_LABEL</type>
<position>68.5,-17.5</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>526</ID>
<type>AA_LABEL</type>
<position>69,-46.5</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>527</ID>
<type>AA_LABEL</type>
<position>155,-5</position>
<gparam>LABEL_TEXT Write MDR input into RAM at MAR address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>528</ID>
<type>AA_LABEL</type>
<position>158.5,-11</position>
<gparam>LABEL_TEXT Write contents of RAM at MAR address to MDR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>529</ID>
<type>AE_REGISTER8</type>
<position>474.5,-20.5</position>
<input>
<ID>IN_0</ID>631 </input>
<input>
<ID>IN_1</ID>630 </input>
<input>
<ID>IN_2</ID>629 </input>
<input>
<ID>IN_3</ID>628 </input>
<input>
<ID>IN_4</ID>627 </input>
<input>
<ID>IN_5</ID>626 </input>
<input>
<ID>IN_6</ID>597 </input>
<input>
<ID>IN_7</ID>640 </input>
<output>
<ID>OUT_0</ID>728 </output>
<output>
<ID>OUT_1</ID>734 </output>
<output>
<ID>OUT_2</ID>520 </output>
<output>
<ID>OUT_3</ID>516 </output>
<output>
<ID>OUT_4</ID>512 </output>
<output>
<ID>OUT_5</ID>508 </output>
<output>
<ID>OUT_6</ID>646 </output>
<output>
<ID>OUT_7</ID>524 </output>
<input>
<ID>clock</ID>642 </input>
<input>
<ID>load</ID>532 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>530</ID>
<type>AE_REGISTER8</type>
<position>128,54</position>
<input>
<ID>IN_0</ID>610 </input>
<input>
<ID>IN_1</ID>611 </input>
<input>
<ID>IN_2</ID>612 </input>
<input>
<ID>IN_3</ID>613 </input>
<input>
<ID>IN_4</ID>614 </input>
<input>
<ID>IN_5</ID>615 </input>
<input>
<ID>IN_6</ID>616 </input>
<input>
<ID>IN_7</ID>617 </input>
<output>
<ID>OUT_0</ID>625 </output>
<output>
<ID>OUT_1</ID>624 </output>
<output>
<ID>OUT_2</ID>623 </output>
<output>
<ID>OUT_3</ID>622 </output>
<output>
<ID>OUT_4</ID>621 </output>
<output>
<ID>OUT_5</ID>620 </output>
<output>
<ID>OUT_6</ID>619 </output>
<output>
<ID>OUT_7</ID>618 </output>
<input>
<ID>clear</ID>609 </input>
<input>
<ID>clock</ID>642 </input>
<input>
<ID>load</ID>608 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>531</ID>
<type>AA_LABEL</type>
<position>120,75.5</position>
<gparam>LABEL_TEXT Global Bus</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>532</ID>
<type>AA_TOGGLE</type>
<position>127,64</position>
<output>
<ID>OUT_0</ID>608 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>533</ID>
<type>AA_LABEL</type>
<position>126.5,67.5</position>
<gparam>LABEL_TEXT Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>534</ID>
<type>AA_TOGGLE</type>
<position>129,45.5</position>
<output>
<ID>OUT_0</ID>609 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>535</ID>
<type>AA_LABEL</type>
<position>129.5,43</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>536</ID>
<type>AA_LABEL</type>
<position>408,45.5</position>
<gparam>LABEL_TEXT SR2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>537</ID>
<type>DA_FROM</type>
<position>108,63</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 7</lparam></gate>
<gate>
<ID>538</ID>
<type>DA_FROM</type>
<position>108.5,59.5</position>
<input>
<ID>IN_0</ID>616 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 6</lparam></gate>
<gate>
<ID>539</ID>
<type>DA_FROM</type>
<position>108,56</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 5</lparam></gate>
<gate>
<ID>540</ID>
<type>DA_FROM</type>
<position>108,53</position>
<input>
<ID>IN_0</ID>614 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 4</lparam></gate>
<gate>
<ID>541</ID>
<type>DA_FROM</type>
<position>108,49.5</position>
<input>
<ID>IN_0</ID>613 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 3</lparam></gate>
<gate>
<ID>542</ID>
<type>DA_FROM</type>
<position>108,46</position>
<input>
<ID>IN_0</ID>612 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 2</lparam></gate>
<gate>
<ID>543</ID>
<type>DA_FROM</type>
<position>108,42.5</position>
<input>
<ID>IN_0</ID>611 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 1</lparam></gate>
<gate>
<ID>544</ID>
<type>DA_FROM</type>
<position>108,39</position>
<input>
<ID>IN_0</ID>610 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 0</lparam></gate>
<gate>
<ID>545</ID>
<type>AE_REGISTER8</type>
<position>476,-44.5</position>
<input>
<ID>IN_0</ID>631 </input>
<input>
<ID>IN_1</ID>630 </input>
<input>
<ID>IN_2</ID>629 </input>
<input>
<ID>IN_3</ID>628 </input>
<input>
<ID>IN_4</ID>627 </input>
<input>
<ID>IN_5</ID>626 </input>
<input>
<ID>IN_6</ID>597 </input>
<input>
<ID>IN_7</ID>640 </input>
<output>
<ID>OUT_0</ID>727 </output>
<output>
<ID>OUT_1</ID>733 </output>
<output>
<ID>OUT_2</ID>521 </output>
<output>
<ID>OUT_3</ID>517 </output>
<output>
<ID>OUT_4</ID>513 </output>
<output>
<ID>OUT_5</ID>509 </output>
<output>
<ID>OUT_6</ID>658 </output>
<output>
<ID>OUT_7</ID>525 </output>
<input>
<ID>clock</ID>642 </input>
<input>
<ID>load</ID>537 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>546</ID>
<type>DE_TO</type>
<position>142.5,64.5</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 7</lparam></gate>
<gate>
<ID>547</ID>
<type>DE_TO</type>
<position>142.5,62</position>
<input>
<ID>IN_0</ID>619 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 6</lparam></gate>
<gate>
<ID>548</ID>
<type>DE_TO</type>
<position>142.5,59.5</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>549</ID>
<type>DE_TO</type>
<position>142.5,56.5</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>550</ID>
<type>DE_TO</type>
<position>142.5,54</position>
<input>
<ID>IN_0</ID>622 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>551</ID>
<type>DE_TO</type>
<position>142.5,50.5</position>
<input>
<ID>IN_0</ID>623 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>552</ID>
<type>DE_TO</type>
<position>142.5,47.5</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>553</ID>
<type>DE_TO</type>
<position>142.5,44.5</position>
<input>
<ID>IN_0</ID>625 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>554</ID>
<type>AE_MUX_4x1</type>
<position>541.5,5.5</position>
<input>
<ID>IN_0</ID>666 </input>
<input>
<ID>IN_1</ID>659 </input>
<input>
<ID>IN_2</ID>658 </input>
<input>
<ID>IN_3</ID>646 </input>
<output>
<ID>OUT</ID>667 </output>
<input>
<ID>SEL_0</ID>595 </input>
<input>
<ID>SEL_1</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>555</ID>
<type>AE_REGISTER8</type>
<position>475.5,-69.5</position>
<input>
<ID>IN_0</ID>631 </input>
<input>
<ID>IN_1</ID>630 </input>
<input>
<ID>IN_2</ID>629 </input>
<input>
<ID>IN_3</ID>628 </input>
<input>
<ID>IN_4</ID>627 </input>
<input>
<ID>IN_5</ID>626 </input>
<input>
<ID>IN_6</ID>597 </input>
<input>
<ID>IN_7</ID>640 </input>
<output>
<ID>OUT_0</ID>670 </output>
<output>
<ID>OUT_1</ID>732 </output>
<output>
<ID>OUT_2</ID>522 </output>
<output>
<ID>OUT_3</ID>518 </output>
<output>
<ID>OUT_4</ID>514 </output>
<output>
<ID>OUT_5</ID>510 </output>
<output>
<ID>OUT_6</ID>659 </output>
<output>
<ID>OUT_7</ID>526 </output>
<input>
<ID>clock</ID>642 </input>
<input>
<ID>load</ID>575 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>556</ID>
<type>AE_MUX_4x1</type>
<position>547.5,-5.5</position>
<input>
<ID>IN_0</ID>666 </input>
<input>
<ID>IN_1</ID>659 </input>
<input>
<ID>IN_2</ID>658 </input>
<input>
<ID>IN_3</ID>646 </input>
<output>
<ID>OUT</ID>668 </output>
<input>
<ID>SEL_0</ID>527 </input>
<input>
<ID>SEL_1</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>557</ID>
<type>AE_REGISTER8</type>
<position>475.5,-94.5</position>
<input>
<ID>IN_0</ID>631 </input>
<input>
<ID>IN_1</ID>630 </input>
<input>
<ID>IN_2</ID>629 </input>
<input>
<ID>IN_3</ID>628 </input>
<input>
<ID>IN_4</ID>627 </input>
<input>
<ID>IN_5</ID>626 </input>
<input>
<ID>IN_6</ID>597 </input>
<input>
<ID>IN_7</ID>640 </input>
<output>
<ID>OUT_0</ID>669 </output>
<output>
<ID>OUT_1</ID>731 </output>
<output>
<ID>OUT_2</ID>523 </output>
<output>
<ID>OUT_3</ID>519 </output>
<output>
<ID>OUT_4</ID>515 </output>
<output>
<ID>OUT_5</ID>511 </output>
<output>
<ID>OUT_6</ID>666 </output>
<output>
<ID>OUT_7</ID>661 </output>
<input>
<ID>clock</ID>642 </input>
<input>
<ID>load</ID>594 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>558</ID>
<type>AA_LABEL</type>
<position>398,-9.5</position>
<gparam>LABEL_TEXT Input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>559</ID>
<type>AA_LABEL</type>
<position>381.5,-79</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>560</ID>
<type>AA_LABEL</type>
<position>408.5,34</position>
<gparam>LABEL_TEXT SR1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>561</ID>
<type>DA_FROM</type>
<position>187,66</position>
<input>
<ID>IN_0</ID>632 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 7</lparam></gate>
<gate>
<ID>562</ID>
<type>DA_FROM</type>
<position>187.5,62.5</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 6</lparam></gate>
<gate>
<ID>563</ID>
<type>DA_FROM</type>
<position>187,59</position>
<input>
<ID>IN_0</ID>634 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>564</ID>
<type>DA_FROM</type>
<position>187,56</position>
<input>
<ID>IN_0</ID>635 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>565</ID>
<type>DA_FROM</type>
<position>187,52.5</position>
<input>
<ID>IN_0</ID>636 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>566</ID>
<type>DA_FROM</type>
<position>187,49</position>
<input>
<ID>IN_0</ID>637 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>567</ID>
<type>DA_FROM</type>
<position>187,45.5</position>
<input>
<ID>IN_0</ID>638 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>568</ID>
<type>DA_FROM</type>
<position>187,42</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>569</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>655,-24</position>
<input>
<ID>IN_0</ID>729 </input>
<input>
<ID>IN_1</ID>735 </input>
<input>
<ID>IN_2</ID>506 </input>
<input>
<ID>IN_3</ID>504 </input>
<input>
<ID>IN_4</ID>502 </input>
<input>
<ID>IN_5</ID>500 </input>
<input>
<ID>IN_6</ID>667 </input>
<input>
<ID>IN_7</ID>596 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>570</ID>
<type>AE_MUX_4x1</type>
<position>608,-119.5</position>
<input>
<ID>IN_0</ID>669 </input>
<input>
<ID>IN_1</ID>670 </input>
<input>
<ID>IN_2</ID>727 </input>
<input>
<ID>IN_3</ID>728 </input>
<output>
<ID>OUT</ID>729 </output>
<input>
<ID>SEL_0</ID>595 </input>
<input>
<ID>SEL_1</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>571</ID>
<type>AE_MUX_4x1</type>
<position>615,-129</position>
<input>
<ID>IN_0</ID>669 </input>
<input>
<ID>IN_1</ID>670 </input>
<input>
<ID>IN_2</ID>727 </input>
<input>
<ID>IN_3</ID>728 </input>
<output>
<ID>OUT</ID>730 </output>
<input>
<ID>SEL_0</ID>527 </input>
<input>
<ID>SEL_1</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>572</ID>
<type>AE_MUX_4x1</type>
<position>585,-78</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>522 </input>
<input>
<ID>IN_2</ID>521 </input>
<input>
<ID>IN_3</ID>520 </input>
<output>
<ID>OUT</ID>506 </output>
<input>
<ID>SEL_0</ID>595 </input>
<input>
<ID>SEL_1</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>573</ID>
<type>AE_MUX_4x1</type>
<position>590.5,-88.5</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>522 </input>
<input>
<ID>IN_2</ID>521 </input>
<input>
<ID>IN_3</ID>520 </input>
<output>
<ID>OUT</ID>507 </output>
<input>
<ID>SEL_0</ID>527 </input>
<input>
<ID>SEL_1</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>574</ID>
<type>AE_MUX_4x1</type>
<position>596,-99</position>
<input>
<ID>IN_0</ID>731 </input>
<input>
<ID>IN_1</ID>732 </input>
<input>
<ID>IN_2</ID>733 </input>
<input>
<ID>IN_3</ID>734 </input>
<output>
<ID>OUT</ID>736 </output>
<input>
<ID>SEL_0</ID>527 </input>
<input>
<ID>SEL_1</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>575</ID>
<type>AE_MUX_4x1</type>
<position>601.5,-109</position>
<input>
<ID>IN_0</ID>731 </input>
<input>
<ID>IN_1</ID>732 </input>
<input>
<ID>IN_2</ID>733 </input>
<input>
<ID>IN_3</ID>734 </input>
<output>
<ID>OUT</ID>735 </output>
<input>
<ID>SEL_0</ID>595 </input>
<input>
<ID>SEL_1</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>576</ID>
<type>DE_TO</type>
<position>177,-27</position>
<input>
<ID>IN_0</ID>600 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 7</lparam></gate>
<gate>
<ID>577</ID>
<type>DE_TO</type>
<position>176,-29.5</position>
<input>
<ID>IN_0</ID>601 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 6</lparam></gate>
<gate>
<ID>578</ID>
<type>DE_TO</type>
<position>176,-32</position>
<input>
<ID>IN_0</ID>602 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 5</lparam></gate>
<gate>
<ID>579</ID>
<type>DA_FROM</type>
<position>210.5,66</position>
<input>
<ID>IN_0</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRsend</lparam></gate>
<gate>
<ID>580</ID>
<type>DE_TO</type>
<position>230.5,-33</position>
<input>
<ID>IN_0</ID>674 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRwrite</lparam></gate>
<gate>
<ID>581</ID>
<type>AA_TOGGLE</type>
<position>221.5,53.5</position>
<output>
<ID>OUT_0</ID>679 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>582</ID>
<type>DE_TO</type>
<position>229,51.5</position>
<input>
<ID>IN_0</ID>679 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 7</lparam></gate>
<gate>
<ID>583</ID>
<type>DE_TO</type>
<position>228,49</position>
<input>
<ID>IN_0</ID>679 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 6</lparam></gate>
<gate>
<ID>584</ID>
<type>DE_TO</type>
<position>228,46.5</position>
<input>
<ID>IN_0</ID>679 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 5</lparam></gate>
<gate>
<ID>585</ID>
<type>DE_TO</type>
<position>228,44</position>
<input>
<ID>IN_0</ID>679 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 4</lparam></gate>
<gate>
<ID>586</ID>
<type>DE_TO</type>
<position>228,41</position>
<input>
<ID>IN_0</ID>678 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 3</lparam></gate>
<gate>
<ID>587</ID>
<type>DE_TO</type>
<position>228.5,38</position>
<input>
<ID>IN_0</ID>677 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 2</lparam></gate>
<gate>
<ID>588</ID>
<type>DE_TO</type>
<position>228.5,35</position>
<input>
<ID>IN_0</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 1</lparam></gate>
<gate>
<ID>589</ID>
<type>DE_TO</type>
<position>228.5,32</position>
<input>
<ID>IN_0</ID>675 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 0</lparam></gate>
<gate>
<ID>590</ID>
<type>DA_FROM</type>
<position>369.5,-9.5</position>
<input>
<ID>IN_0</ID>683 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID REGin</lparam></gate>
<gate>
<ID>591</ID>
<type>DE_TO</type>
<position>233,-30</position>
<input>
<ID>IN_0</ID>684 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID REGin</lparam></gate>
<gate>
<ID>592</ID>
<type>DD_KEYPAD_HEX</type>
<position>271,-144</position>
<output>
<ID>OUT_0</ID>697 </output>
<output>
<ID>OUT_1</ID>696 </output>
<output>
<ID>OUT_2</ID>695 </output>
<output>
<ID>OUT_3</ID>694 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>593</ID>
<type>DD_KEYPAD_HEX</type>
<position>271,-159</position>
<output>
<ID>OUT_0</ID>693 </output>
<output>
<ID>OUT_1</ID>692 </output>
<output>
<ID>OUT_2</ID>691 </output>
<output>
<ID>OUT_3</ID>690 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>594</ID>
<type>DD_KEYPAD_HEX</type>
<position>271,-173.5</position>
<output>
<ID>OUT_0</ID>701 </output>
<output>
<ID>OUT_1</ID>700 </output>
<output>
<ID>OUT_2</ID>699 </output>
<output>
<ID>OUT_3</ID>698 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>595</ID>
<type>AA_AND2</type>
<position>310,-161</position>
<input>
<ID>IN_0</ID>686 </input>
<input>
<ID>IN_1</ID>690 </input>
<output>
<ID>OUT</ID>710 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>596</ID>
<type>AA_AND2</type>
<position>310,-166.5</position>
<input>
<ID>IN_0</ID>687 </input>
<input>
<ID>IN_1</ID>691 </input>
<output>
<ID>OUT</ID>711 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>597</ID>
<type>AA_AND2</type>
<position>310,-172</position>
<input>
<ID>IN_0</ID>688 </input>
<input>
<ID>IN_1</ID>692 </input>
<output>
<ID>OUT</ID>712 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>598</ID>
<type>AA_AND2</type>
<position>310,-177.5</position>
<input>
<ID>IN_0</ID>689 </input>
<input>
<ID>IN_1</ID>693 </input>
<output>
<ID>OUT</ID>713 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>599</ID>
<type>AA_AND2</type>
<position>310,-183</position>
<input>
<ID>IN_0</ID>694 </input>
<input>
<ID>IN_1</ID>698 </input>
<output>
<ID>OUT</ID>714 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>600</ID>
<type>AA_AND2</type>
<position>310,-188.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>699 </input>
<output>
<ID>OUT</ID>715 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>601</ID>
<type>AA_AND2</type>
<position>310,-193.5</position>
<input>
<ID>IN_0</ID>696 </input>
<input>
<ID>IN_1</ID>700 </input>
<output>
<ID>OUT</ID>716 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>602</ID>
<type>AA_AND2</type>
<position>310,-199</position>
<input>
<ID>IN_0</ID>697 </input>
<input>
<ID>IN_1</ID>701 </input>
<output>
<ID>OUT</ID>717 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>603</ID>
<type>AA_MUX_2x1</type>
<position>337.5,-142</position>
<input>
<ID>IN_0</ID>709 </input>
<input>
<ID>IN_1</ID>717 </input>
<output>
<ID>OUT</ID>719 </output>
<input>
<ID>SEL_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>604</ID>
<type>AA_MUX_2x1</type>
<position>337.5,-147.5</position>
<input>
<ID>IN_0</ID>708 </input>
<input>
<ID>IN_1</ID>716 </input>
<output>
<ID>OUT</ID>720 </output>
<input>
<ID>SEL_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>605</ID>
<type>AA_MUX_2x1</type>
<position>337.5,-153</position>
<input>
<ID>IN_0</ID>707 </input>
<input>
<ID>IN_1</ID>715 </input>
<output>
<ID>OUT</ID>721 </output>
<input>
<ID>SEL_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>606</ID>
<type>AA_MUX_2x1</type>
<position>337.5,-158</position>
<input>
<ID>IN_0</ID>706 </input>
<input>
<ID>IN_1</ID>714 </input>
<output>
<ID>OUT</ID>722 </output>
<input>
<ID>SEL_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>607</ID>
<type>AA_MUX_2x1</type>
<position>337.5,-168.5</position>
<input>
<ID>IN_0</ID>705 </input>
<input>
<ID>IN_1</ID>713 </input>
<output>
<ID>OUT</ID>723 </output>
<input>
<ID>SEL_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>608</ID>
<type>AA_MUX_2x1</type>
<position>337.5,-173.5</position>
<input>
<ID>IN_0</ID>704 </input>
<input>
<ID>IN_1</ID>712 </input>
<output>
<ID>OUT</ID>724 </output>
<input>
<ID>SEL_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>609</ID>
<type>AA_MUX_2x1</type>
<position>337.5,-178.5</position>
<input>
<ID>IN_0</ID>703 </input>
<input>
<ID>IN_1</ID>711 </input>
<output>
<ID>OUT</ID>725 </output>
<input>
<ID>SEL_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>610</ID>
<type>AA_MUX_2x1</type>
<position>337.5,-183.5</position>
<input>
<ID>IN_0</ID>702 </input>
<input>
<ID>IN_1</ID>710 </input>
<output>
<ID>OUT</ID>726 </output>
<input>
<ID>SEL_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>611</ID>
<type>AA_TOGGLE</type>
<position>341,-128.5</position>
<output>
<ID>OUT_0</ID>718 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>612</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>368,-163.5</position>
<input>
<ID>IN_0</ID>726 </input>
<input>
<ID>IN_1</ID>725 </input>
<input>
<ID>IN_2</ID>724 </input>
<input>
<ID>IN_3</ID>723 </input>
<input>
<ID>IN_4</ID>722 </input>
<input>
<ID>IN_5</ID>721 </input>
<input>
<ID>IN_6</ID>720 </input>
<input>
<ID>IN_7</ID>719 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 136</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>613</ID>
<type>AA_LABEL</type>
<position>260.5,-137</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>614</ID>
<type>AA_LABEL</type>
<position>261.5,-165.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>615</ID>
<type>AA_LABEL</type>
<position>354,-128</position>
<gparam>LABEL_TEXT Control Signal</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>616</ID>
<type>AE_FULLADDER_4BIT</type>
<position>310.5,-134.5</position>
<input>
<ID>IN_0</ID>697 </input>
<input>
<ID>IN_1</ID>696 </input>
<input>
<ID>IN_2</ID>695 </input>
<input>
<ID>IN_3</ID>694 </input>
<input>
<ID>IN_B_0</ID>701 </input>
<input>
<ID>IN_B_1</ID>700 </input>
<input>
<ID>IN_B_2</ID>699 </input>
<input>
<ID>IN_B_3</ID>698 </input>
<output>
<ID>OUT_0</ID>702 </output>
<output>
<ID>OUT_1</ID>703 </output>
<output>
<ID>OUT_2</ID>704 </output>
<output>
<ID>OUT_3</ID>705 </output>
<output>
<ID>carry_out</ID>685 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>617</ID>
<type>AE_FULLADDER_4BIT</type>
<position>310.5,-150.5</position>
<input>
<ID>IN_0</ID>689 </input>
<input>
<ID>IN_1</ID>688 </input>
<input>
<ID>IN_2</ID>687 </input>
<input>
<ID>IN_3</ID>686 </input>
<input>
<ID>IN_B_0</ID>693 </input>
<input>
<ID>IN_B_1</ID>692 </input>
<input>
<ID>IN_B_2</ID>691 </input>
<input>
<ID>IN_B_3</ID>690 </input>
<output>
<ID>OUT_0</ID>706 </output>
<output>
<ID>OUT_1</ID>707 </output>
<output>
<ID>OUT_2</ID>708 </output>
<output>
<ID>OUT_3</ID>709 </output>
<input>
<ID>carry_in</ID>685 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>618</ID>
<type>DD_KEYPAD_HEX</type>
<position>271,-130.5</position>
<output>
<ID>OUT_0</ID>689 </output>
<output>
<ID>OUT_1</ID>688 </output>
<output>
<ID>OUT_2</ID>687 </output>
<output>
<ID>OUT_3</ID>686 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>619</ID>
<type>DE_TO</type>
<position>176,-34.5</position>
<input>
<ID>IN_0</ID>603 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 4</lparam></gate>
<gate>
<ID>620</ID>
<type>DE_TO</type>
<position>176,-37.5</position>
<input>
<ID>IN_0</ID>604 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 3</lparam></gate>
<gate>
<ID>621</ID>
<type>DE_TO</type>
<position>176.5,-40.5</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 2</lparam></gate>
<gate>
<ID>622</ID>
<type>DE_TO</type>
<position>176.5,-43.5</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 1</lparam></gate>
<gate>
<ID>623</ID>
<type>DE_TO</type>
<position>176.5,-46.5</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 0</lparam></gate>
<gate>
<ID>624</ID>
<type>BB_CLOCK</type>
<position>172,24.5</position>
<output>
<ID>CLK</ID>642 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>625</ID>
<type>DA_FROM</type>
<position>90,-33.5</position>
<input>
<ID>IN_0</ID>593 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 7</lparam></gate>
<gate>
<ID>626</ID>
<type>DA_FROM</type>
<position>90,-40.5</position>
<input>
<ID>IN_0</ID>644 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>627</ID>
<type>DA_FROM</type>
<position>90,-43.5</position>
<input>
<ID>IN_0</ID>645 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>628</ID>
<type>DA_FROM</type>
<position>90,-47</position>
<input>
<ID>IN_0</ID>648 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>629</ID>
<type>DA_FROM</type>
<position>90,-50.5</position>
<input>
<ID>IN_0</ID>647 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>630</ID>
<type>DA_FROM</type>
<position>90,-54</position>
<input>
<ID>IN_0</ID>598 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>631</ID>
<type>DA_FROM</type>
<position>90,-57.5</position>
<input>
<ID>IN_0</ID>599 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>632</ID>
<type>DA_FROM</type>
<position>89.5,-37.5</position>
<input>
<ID>IN_0</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 6</lparam></gate>
<gate>
<ID>633</ID>
<type>DE_TO</type>
<position>337.5,42</position>
<input>
<ID>IN_0</ID>657 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 7</lparam></gate>
<gate>
<ID>634</ID>
<type>DE_TO</type>
<position>336.5,39.5</position>
<input>
<ID>IN_0</ID>656 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 6</lparam></gate>
<gate>
<ID>635</ID>
<type>DE_TO</type>
<position>336.5,37</position>
<input>
<ID>IN_0</ID>655 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 5</lparam></gate>
<gate>
<ID>636</ID>
<type>DE_TO</type>
<position>336.5,34.5</position>
<input>
<ID>IN_0</ID>654 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 4</lparam></gate>
<gate>
<ID>637</ID>
<type>DE_TO</type>
<position>336.5,31.5</position>
<input>
<ID>IN_0</ID>653 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 3</lparam></gate>
<gate>
<ID>638</ID>
<type>DE_TO</type>
<position>337,28.5</position>
<input>
<ID>IN_0</ID>652 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 2</lparam></gate>
<gate>
<ID>639</ID>
<type>DE_TO</type>
<position>337,25.5</position>
<input>
<ID>IN_0</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 1</lparam></gate>
<gate>
<ID>640</ID>
<type>DE_TO</type>
<position>337,22.5</position>
<input>
<ID>IN_0</ID>649 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 0</lparam></gate>
<gate>
<ID>641</ID>
<type>AE_MUX_4x1</type>
<position>553.5,-15.5</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>510 </input>
<input>
<ID>IN_2</ID>509 </input>
<input>
<ID>IN_3</ID>508 </input>
<output>
<ID>OUT</ID>500 </output>
<input>
<ID>SEL_0</ID>595 </input>
<input>
<ID>SEL_1</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>642</ID>
<type>AA_LABEL</type>
<position>344.5,49.5</position>
<gparam>LABEL_TEXT Send PC to Bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>643</ID>
<type>AE_MUX_4x1</type>
<position>559,-26.5</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>510 </input>
<input>
<ID>IN_2</ID>509 </input>
<input>
<ID>IN_3</ID>508 </input>
<output>
<ID>OUT</ID>501 </output>
<input>
<ID>SEL_0</ID>527 </input>
<input>
<ID>SEL_1</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>644</ID>
<type>BI_ROM_12x16</type>
<position>228.5,-8.5</position>
<input>
<ID>ADDRESS_0</ID>680 </input>
<input>
<ID>ADDRESS_1</ID>681 </input>
<input>
<ID>ADDRESS_2</ID>682 </input>
<input>
<ID>ADDRESS_3</ID>660 </input>
<input>
<ID>ADDRESS_4</ID>671 </input>
<input>
<ID>ADDRESS_5</ID>672 </input>
<output>
<ID>DATA_OUT_0</ID>680 </output>
<output>
<ID>DATA_OUT_1</ID>681 </output>
<output>
<ID>DATA_OUT_10</ID>536 </output>
<output>
<ID>DATA_OUT_11</ID>737 </output>
<output>
<ID>DATA_OUT_12</ID>664 </output>
<output>
<ID>DATA_OUT_13</ID>665 </output>
<output>
<ID>DATA_OUT_14</ID>663 </output>
<output>
<ID>DATA_OUT_15</ID>662 </output>
<output>
<ID>DATA_OUT_2</ID>682 </output>
<output>
<ID>DATA_OUT_8</ID>684 </output>
<output>
<ID>DATA_OUT_9</ID>674 </output>
<input>
<ID>ENABLE_0</ID>742 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam></gate>
<gate>
<ID>645</ID>
<type>AE_MUX_4x1</type>
<position>528,23.5</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>526 </input>
<input>
<ID>IN_2</ID>525 </input>
<input>
<ID>IN_3</ID>524 </input>
<output>
<ID>OUT</ID>596 </output>
<input>
<ID>SEL_0</ID>595 </input>
<input>
<ID>SEL_1</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>646</ID>
<type>AE_MUX_4x1</type>
<position>564,-37</position>
<input>
<ID>IN_0</ID>515 </input>
<input>
<ID>IN_1</ID>514 </input>
<input>
<ID>IN_2</ID>513 </input>
<input>
<ID>IN_3</ID>512 </input>
<output>
<ID>OUT</ID>502 </output>
<input>
<ID>SEL_0</ID>595 </input>
<input>
<ID>SEL_1</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>647</ID>
<type>AA_LABEL</type>
<position>386.5,-94</position>
<gparam>LABEL_TEXT DR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>648</ID>
<type>AE_MUX_4x1</type>
<position>569.5,-47</position>
<input>
<ID>IN_0</ID>515 </input>
<input>
<ID>IN_1</ID>514 </input>
<input>
<ID>IN_2</ID>513 </input>
<input>
<ID>IN_3</ID>512 </input>
<output>
<ID>OUT</ID>503 </output>
<input>
<ID>SEL_0</ID>527 </input>
<input>
<ID>SEL_1</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>649</ID>
<type>AE_MUX_4x1</type>
<position>575,-57.5</position>
<input>
<ID>IN_0</ID>519 </input>
<input>
<ID>IN_1</ID>518 </input>
<input>
<ID>IN_2</ID>517 </input>
<input>
<ID>IN_3</ID>516 </input>
<output>
<ID>OUT</ID>504 </output>
<input>
<ID>SEL_0</ID>595 </input>
<input>
<ID>SEL_1</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>650</ID>
<type>AE_MUX_4x1</type>
<position>580.5,-68</position>
<input>
<ID>IN_0</ID>519 </input>
<input>
<ID>IN_1</ID>518 </input>
<input>
<ID>IN_2</ID>517 </input>
<input>
<ID>IN_3</ID>516 </input>
<output>
<ID>OUT</ID>505 </output>
<input>
<ID>SEL_0</ID>527 </input>
<input>
<ID>SEL_1</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>651</ID>
<type>AA_TOGGLE</type>
<position>391,-93.5</position>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>652</ID>
<type>DE_TO</type>
<position>223.5,-54</position>
<input>
<ID>IN_0</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID sendPC</lparam></gate>
<gate>
<ID>653</ID>
<type>DA_FROM</type>
<position>326.5,53</position>
<input>
<ID>IN_0</ID>651 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID sendPC</lparam></gate>
<gate>
<ID>654</ID>
<type>DA_FROM</type>
<position>90.5,-5</position>
<input>
<ID>IN_0</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 7</lparam></gate>
<gate>
<ID>655</ID>
<type>DA_FROM</type>
<position>90.5,-12</position>
<input>
<ID>IN_0</ID>550 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>656</ID>
<type>DA_FROM</type>
<position>90.5,-15</position>
<input>
<ID>IN_0</ID>551 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>657</ID>
<type>DA_FROM</type>
<position>90.5,-18.5</position>
<input>
<ID>IN_0</ID>552 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>658</ID>
<type>DA_FROM</type>
<position>90.5,-22</position>
<input>
<ID>IN_0</ID>553 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>659</ID>
<type>DA_FROM</type>
<position>90.5,-25.5</position>
<input>
<ID>IN_0</ID>554 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>660</ID>
<type>DA_FROM</type>
<position>90.5,-29</position>
<input>
<ID>IN_0</ID>555 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>661</ID>
<type>DA_FROM</type>
<position>90.5,-9</position>
<input>
<ID>IN_0</ID>549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 6</lparam></gate>
<gate>
<ID>662</ID>
<type>BA_DECODER_2x4</type>
<position>401.5,-87</position>
<input>
<ID>ENABLE</ID>683 </input>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>530 </input>
<output>
<ID>OUT_0</ID>594 </output>
<output>
<ID>OUT_1</ID>575 </output>
<output>
<ID>OUT_2</ID>537 </output>
<output>
<ID>OUT_3</ID>532 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>663</ID>
<type>DA_FROM</type>
<position>128.5,-6</position>
<input>
<ID>IN_0</ID>592 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRwrite</lparam></gate>
<gate>
<ID>664</ID>
<type>AE_MUX_4x1</type>
<position>534,14</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>526 </input>
<input>
<ID>IN_2</ID>525 </input>
<input>
<ID>IN_3</ID>524 </input>
<output>
<ID>OUT</ID>641 </output>
<input>
<ID>SEL_0</ID>527 </input>
<input>
<ID>SEL_1</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>665</ID>
<type>DA_FROM</type>
<position>140,-13.5</position>
<input>
<ID>IN_0</ID>743 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID MAR</lparam></gate>
<gate>
<ID>666</ID>
<type>DE_TO</type>
<position>224,-50.5</position>
<input>
<ID>IN_0</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR</lparam></gate>
<gate>
<ID>667</ID>
<type>AA_LABEL</type>
<position>307,-116</position>
<gparam>LABEL_TEXT ALU</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>323</ID>
<type>DE_TO</type>
<position>225.5,-46.5</position>
<input>
<ID>IN_0</ID>665 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRload</lparam></gate>
<gate>
<ID>324</ID>
<type>DE_TO</type>
<position>226,-42</position>
<input>
<ID>IN_0</ID>664 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRsend</lparam></gate>
<gate>
<ID>325</ID>
<type>DA_FROM</type>
<position>188.5,70.5</position>
<input>
<ID>IN_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRrecieve</lparam></gate>
<gate>
<ID>326</ID>
<type>DD_KEYPAD_HEX</type>
<position>77,-106</position>
<output>
<ID>OUT_0</ID>424 </output>
<output>
<ID>OUT_1</ID>423 </output>
<output>
<ID>OUT_2</ID>422 </output>
<output>
<ID>OUT_3</ID>421 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>327</ID>
<type>DE_TO</type>
<position>86,-101.5</position>
<input>
<ID>IN_0</ID>421 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 0</lparam></gate>
<gate>
<ID>328</ID>
<type>DE_TO</type>
<position>86,-104.5</position>
<input>
<ID>IN_0</ID>422 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 1</lparam></gate>
<gate>
<ID>329</ID>
<type>DE_TO</type>
<position>86,-107.5</position>
<input>
<ID>IN_0</ID>423 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 2</lparam></gate>
<gate>
<ID>330</ID>
<type>DE_TO</type>
<position>86,-110.5</position>
<input>
<ID>IN_0</ID>424 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 3</lparam></gate>
<gate>
<ID>331</ID>
<type>DE_TO</type>
<position>86,-113.5</position>
<input>
<ID>IN_0</ID>424 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 4</lparam></gate>
<gate>
<ID>332</ID>
<type>DE_TO</type>
<position>86,-116.5</position>
<input>
<ID>IN_0</ID>424 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 5</lparam></gate>
<gate>
<ID>333</ID>
<type>DE_TO</type>
<position>86,-119.5</position>
<input>
<ID>IN_0</ID>424 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 6</lparam></gate>
<gate>
<ID>334</ID>
<type>DE_TO</type>
<position>86,-122.5</position>
<input>
<ID>IN_0</ID>424 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 7</lparam></gate>
<gate>
<ID>335</ID>
<type>AA_TOGGLE</type>
<position>211,-149</position>
<output>
<ID>OUT_0</ID>462 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_FULLADDER_4BIT</type>
<position>186,-118</position>
<input>
<ID>IN_0</ID>454 </input>
<input>
<ID>IN_1</ID>455 </input>
<input>
<ID>IN_2</ID>456 </input>
<input>
<ID>IN_3</ID>457 </input>
<input>
<ID>IN_B_0</ID>453 </input>
<input>
<ID>IN_B_1</ID>452 </input>
<input>
<ID>IN_B_2</ID>451 </input>
<input>
<ID>IN_B_3</ID>450 </input>
<output>
<ID>OUT_0</ID>460 </output>
<output>
<ID>OUT_1</ID>459 </output>
<output>
<ID>OUT_2</ID>458 </output>
<output>
<ID>OUT_3</ID>466 </output>
<output>
<ID>carry_out</ID>483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>337</ID>
<type>AE_FULLADDER_4BIT</type>
<position>132,-118</position>
<input>
<ID>IN_0</ID>425 </input>
<input>
<ID>IN_1</ID>426 </input>
<input>
<ID>IN_2</ID>427 </input>
<input>
<ID>IN_3</ID>428 </input>
<input>
<ID>IN_B_0</ID>429 </input>
<input>
<ID>IN_B_1</ID>430 </input>
<input>
<ID>IN_B_2</ID>431 </input>
<input>
<ID>IN_B_3</ID>448 </input>
<output>
<ID>OUT_0</ID>472 </output>
<output>
<ID>OUT_1</ID>474 </output>
<output>
<ID>OUT_2</ID>475 </output>
<output>
<ID>OUT_3</ID>476 </output>
<input>
<ID>carry_in</ID>483 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>361</ID>
<type>DE_TO</type>
<position>227,-38</position>
<input>
<ID>IN_0</ID>737 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRrecieve</lparam></gate>
<gate>
<ID>373</ID>
<type>AA_MUX_2x1</type>
<position>178.5,-134</position>
<input>
<ID>IN_0</ID>467 </input>
<input>
<ID>IN_1</ID>458 </input>
<output>
<ID>OUT</ID>468 </output>
<input>
<ID>SEL_0</ID>462 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>387</ID>
<type>AA_MUX_2x1</type>
<position>151.5,-140</position>
<input>
<ID>IN_0</ID>471 </input>
<input>
<ID>IN_1</ID>472 </input>
<output>
<ID>OUT</ID>473 </output>
<input>
<ID>SEL_0</ID>462 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>421</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-103,83,-103</points>
<connection>
<GID>326</GID>
<name>OUT_3</name></connection>
<intersection>83 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83,-103,83,-101.5</points>
<intersection>-103 1</intersection>
<intersection>-101.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>83,-101.5,84,-101.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>83 3</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-105,83,-104.5</points>
<intersection>-105 2</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-104.5,84,-104.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-105,83,-105</points>
<connection>
<GID>326</GID>
<name>OUT_2</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-107.5,83,-107</points>
<intersection>-107.5 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-107.5,84,-107.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-107,83,-107</points>
<connection>
<GID>326</GID>
<name>OUT_1</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-109,83,-109</points>
<connection>
<GID>326</GID>
<name>OUT_0</name></connection>
<intersection>83 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83,-122.5,83,-109</points>
<intersection>-122.5 8</intersection>
<intersection>-119.5 9</intersection>
<intersection>-116.5 10</intersection>
<intersection>-113.5 11</intersection>
<intersection>-110.5 12</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>83,-122.5,84,-122.5</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>83 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>83,-119.5,84,-119.5</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>83 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>83,-116.5,84,-116.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>83 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>83,-113.5,84,-113.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>83 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>83,-110.5,84,-110.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>83 3</intersection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-114,130,-111</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>-111 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,-111,130.5,-111</points>
<intersection>130 0</intersection>
<intersection>130.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>130.5,-111,130.5,-110</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>-111 3</intersection></vsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-114,129,-111</points>
<connection>
<GID>337</GID>
<name>IN_1</name></connection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-111,129,-111</points>
<intersection>127.5 4</intersection>
<intersection>129 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127.5,-111,127.5,-110</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>-111 2</intersection></vsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>124.5,-112,128,-112</points>
<intersection>124.5 4</intersection>
<intersection>128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128,-114,128,-112</points>
<connection>
<GID>337</GID>
<name>IN_2</name></connection>
<intersection>-112 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>124.5,-112,124.5,-110</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>-112 2</intersection></vsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>121.5,-113,127,-113</points>
<intersection>121.5 5</intersection>
<intersection>127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127,-114,127,-113</points>
<connection>
<GID>337</GID>
<name>IN_3</name></connection>
<intersection>-113 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>121.5,-113,121.5,-110</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>-113 2</intersection></vsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>142.5,-113,142.5,-110</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>137,-113,142.5,-113</points>
<intersection>137 3</intersection>
<intersection>142.5 1</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>137,-114,137,-113</points>
<connection>
<GID>337</GID>
<name>IN_B_0</name></connection>
<intersection>-113 2</intersection></vsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-114,136,-112</points>
<connection>
<GID>337</GID>
<name>IN_B_1</name></connection>
<intersection>-112 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>139.5,-112,139.5,-110</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>136,-112,139.5,-112</points>
<intersection>136 0</intersection>
<intersection>139.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-111,136.5,-110</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>-111 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>135,-114,135,-111</points>
<connection>
<GID>337</GID>
<name>IN_B_2</name></connection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>135,-111,136.5,-111</points>
<intersection>135 1</intersection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>134,-114,134,-111</points>
<connection>
<GID>337</GID>
<name>IN_B_3</name></connection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>133.5,-111,134,-111</points>
<intersection>133.5 4</intersection>
<intersection>134 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>133.5,-111,133.5,-110</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>-111 2</intersection></vsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-114,188,-111</points>
<connection>
<GID>336</GID>
<name>IN_B_3</name></connection>
<intersection>-111 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>187.5,-111,188,-111</points>
<intersection>187.5 5</intersection>
<intersection>188 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>187.5,-111,187.5,-110</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>-111 3</intersection></vsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-111,190.5,-110</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>-111 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>189,-114,189,-111</points>
<connection>
<GID>336</GID>
<name>IN_B_2</name></connection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>189,-111,190.5,-111</points>
<intersection>189 1</intersection>
<intersection>190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-114,190,-112</points>
<connection>
<GID>336</GID>
<name>IN_B_1</name></connection>
<intersection>-112 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>193.5,-112,193.5,-110</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>190,-112,193.5,-112</points>
<intersection>190 0</intersection>
<intersection>193.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-114,191,-113</points>
<connection>
<GID>336</GID>
<name>IN_B_0</name></connection>
<intersection>-113 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>196.5,-113,196.5,-110</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>191,-113,196.5,-113</points>
<intersection>191 0</intersection>
<intersection>196.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-114,184,-111</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>-111 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>184.5,-111,184.5,-110</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>184,-111,184.5,-111</points>
<intersection>184 0</intersection>
<intersection>184.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-114,183,-111</points>
<connection>
<GID>336</GID>
<name>IN_1</name></connection>
<intersection>-111 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>181.5,-111,181.5,-110</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>181.5,-111,183,-111</points>
<intersection>181.5 1</intersection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,-114,182,-112</points>
<connection>
<GID>336</GID>
<name>IN_2</name></connection>
<intersection>-112 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>178.5,-112,178.5,-110</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-112,182,-112</points>
<intersection>178.5 1</intersection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>175.5,-113,175.5,-110</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>175.5,-113,181,-113</points>
<intersection>175.5 1</intersection>
<intersection>181 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>181,-114,181,-113</points>
<connection>
<GID>336</GID>
<name>IN_3</name></connection>
<intersection>-113 2</intersection></vsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>179.5,-124,185.5,-124</points>
<intersection>179.5 13</intersection>
<intersection>185.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>185.5,-124,185.5,-122</points>
<connection>
<GID>336</GID>
<name>OUT_2</name></connection>
<intersection>-124 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>179.5,-132,179.5,-124</points>
<connection>
<GID>373</GID>
<name>IN_1</name></connection>
<intersection>-124 11</intersection></vsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,-129,192.5,-124</points>
<connection>
<GID>403</GID>
<name>IN_1</name></connection>
<intersection>-124 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>186.5,-124,192.5,-124</points>
<intersection>186.5 17</intersection>
<intersection>192.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>186.5,-124,186.5,-122</points>
<connection>
<GID>336</GID>
<name>OUT_1</name></connection>
<intersection>-124 16</intersection></vsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-123,187.5,-122</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>187.5,-123,206.5,-123</points>
<intersection>187.5 0</intersection>
<intersection>206.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>206.5,-126,206.5,-123</points>
<connection>
<GID>394</GID>
<name>IN_1</name></connection>
<intersection>-123 2</intersection></vsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203.5,-125,204.5,-125</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>204.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>204.5,-126,204.5,-125</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>-125 1</intersection></vsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-149,209,-149</points>
<connection>
<GID>396</GID>
<name>SEL_0</name></connection>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>126 34</intersection>
<intersection>139.5 32</intersection>
<intersection>152.5 28</intersection>
<intersection>166.5 22</intersection>
<intersection>180 13</intersection>
<intersection>193 8</intersection>
<intersection>207 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>207,-149,207,-128</points>
<intersection>-149 1</intersection>
<intersection>-128 38</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>193,-149,193,-131</points>
<intersection>-149 1</intersection>
<intersection>-131 42</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>180,-149,180,-134</points>
<intersection>-149 1</intersection>
<intersection>-134 36</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>166.5,-149,166.5,-137</points>
<intersection>-149 1</intersection>
<intersection>-137 40</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>152.5,-149,152.5,-140</points>
<intersection>-149 1</intersection>
<intersection>-140 44</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>139.5,-149,139.5,-143</points>
<intersection>-149 1</intersection>
<intersection>-143 37</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>126,-149,126,-146</points>
<intersection>-149 1</intersection>
<intersection>-146 41</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>180,-134,181,-134</points>
<connection>
<GID>373</GID>
<name>SEL_0</name></connection>
<intersection>180 13</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>139.5,-143,140.5,-143</points>
<connection>
<GID>391</GID>
<name>SEL_0</name></connection>
<intersection>139.5 32</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>207,-128,208,-128</points>
<connection>
<GID>394</GID>
<name>SEL_0</name></connection>
<intersection>207 4</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>166.5,-137,167.5,-137</points>
<connection>
<GID>397</GID>
<name>SEL_0</name></connection>
<intersection>166.5 22</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>126,-146,127,-146</points>
<connection>
<GID>402</GID>
<name>SEL_0</name></connection>
<intersection>126 34</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>193,-131,194,-131</points>
<connection>
<GID>403</GID>
<name>SEL_0</name></connection>
<intersection>193 8</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>152.5,-140,154,-140</points>
<connection>
<GID>387</GID>
<name>SEL_0</name></connection>
<intersection>152.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-152,205.5,-130</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<connection>
<GID>394</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-129,190.5,-126</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>-126 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>190,-126,190.5,-126</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-152,191.5,-133</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<connection>
<GID>403</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-135,166,-123</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>-123 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>184.5,-123,184.5,-122</points>
<connection>
<GID>336</GID>
<name>OUT_3</name></connection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>166,-123,184.5,-123</points>
<intersection>166 0</intersection>
<intersection>184.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177.5,-132,177.5,-125</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>-125 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>176.5,-125,177.5,-125</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>177.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-152,178.5,-136</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<connection>
<GID>373</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-152,165,-139</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<connection>
<GID>397</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164,-135,164,-124</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>-124 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>163,-124,164,-124</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>164 0</intersection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-138,150.5,-125</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>-125 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>149.5,-125,150.5,-125</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-138,152.5,-123</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<intersection>-123 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>133.5,-123,133.5,-122</points>
<connection>
<GID>337</GID>
<name>OUT_0</name></connection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>133.5,-123,152.5,-123</points>
<intersection>133.5 1</intersection>
<intersection>152.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-152,151.5,-142</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<connection>
<GID>387</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-141,139,-124</points>
<connection>
<GID>391</GID>
<name>IN_1</name></connection>
<intersection>-124 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>132.5,-124,139,-124</points>
<intersection>132.5 4</intersection>
<intersection>139 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>132.5,-124,132.5,-122</points>
<connection>
<GID>337</GID>
<name>OUT_1</name></connection>
<intersection>-124 3</intersection></vsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-124,131.5,-122</points>
<connection>
<GID>337</GID>
<name>OUT_2</name></connection>
<intersection>-124 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>125.5,-144,125.5,-124</points>
<connection>
<GID>402</GID>
<name>IN_1</name></connection>
<intersection>-124 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-124,131.5,-124</points>
<intersection>125.5 1</intersection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-123,130.5,-122</points>
<connection>
<GID>337</GID>
<name>OUT_3</name></connection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>112,-123,130.5,-123</points>
<intersection>112 3</intersection>
<intersection>130.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>112,-147,112,-123</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<intersection>-123 2</intersection></vsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-141,137,-126</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>-126 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>136,-126,137,-126</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-144,123.5,-125</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>-125 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>122.5,-125,123.5,-125</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-147,110,-124</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>-124 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>109,-124,110,-124</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-152,138,-145</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<connection>
<GID>391</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-152,124.5,-148</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<connection>
<GID>402</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>111,-152,111,-151</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<connection>
<GID>396</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140,-117,178,-117</points>
<connection>
<GID>337</GID>
<name>carry_in</name></connection>
<connection>
<GID>336</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>375,-55.5,375,-40</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>-55.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>367.5,-55.5,375,-55.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>375 11</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373.5,-47.5,373.5,-39</points>
<intersection>-47.5 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>373.5,-39,375,-39</points>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<intersection>373.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>368,-47.5,373.5,-47.5</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>373.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-42.5,372,-38</points>
<intersection>-42.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>365.5,-42.5,372,-42.5</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>372 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372,-38,375,-38</points>
<connection>
<GID>450</GID>
<name>IN_2</name></connection>
<intersection>372 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>363.5,-37,375,-37</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<connection>
<GID>450</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,-36,366.5,-33</points>
<intersection>-36 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>366.5,-36,375,-36</points>
<connection>
<GID>450</GID>
<name>IN_4</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>346.5,-33,366.5,-33</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>366.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368,-35,368,-31</points>
<intersection>-35 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>368,-35,375,-35</points>
<connection>
<GID>450</GID>
<name>IN_5</name></connection>
<intersection>368 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347.5,-31,368,-31</points>
<intersection>347.5 3</intersection>
<intersection>368 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>347.5,-31,347.5,-27.5</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>371,-34,371,-23.5</points>
<intersection>-34 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>371,-34,375,-34</points>
<connection>
<GID>450</GID>
<name>IN_6</name></connection>
<intersection>371 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347,-23.5,371,-23.5</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>371 0</intersection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373.5,-33,373.5,-19.5</points>
<intersection>-33 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>373.5,-33,375,-33</points>
<connection>
<GID>450</GID>
<name>IN_7</name></connection>
<intersection>373.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347,-19.5,373.5,-19.5</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>373.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>145,-36.5,145,-36</points>
<connection>
<GID>470</GID>
<name>clear</name></connection>
<intersection>-36.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>143,-36.5,145,-36.5</points>
<intersection>143 11</intersection>
<intersection>145 4</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>143,-37.5,143,-36.5</points>
<connection>
<GID>488</GID>
<name>OUT_0</name></connection>
<intersection>-36.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-25.5,157.5,-23</points>
<connection>
<GID>495</GID>
<name>ENABLE_0</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-23,158.5,-23</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>148,-27,155.5,-27</points>
<connection>
<GID>470</GID>
<name>OUT_7</name></connection>
<connection>
<GID>495</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>148,-28,155.5,-28</points>
<connection>
<GID>470</GID>
<name>OUT_6</name></connection>
<connection>
<GID>495</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>148,-29,155.5,-29</points>
<connection>
<GID>470</GID>
<name>OUT_5</name></connection>
<connection>
<GID>495</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>148,-30,155.5,-30</points>
<connection>
<GID>470</GID>
<name>OUT_4</name></connection>
<connection>
<GID>495</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>148,-31,155.5,-31</points>
<connection>
<GID>470</GID>
<name>OUT_3</name></connection>
<connection>
<GID>495</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>148,-32,155.5,-32</points>
<connection>
<GID>470</GID>
<name>OUT_2</name></connection>
<connection>
<GID>495</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>603,-22,603,-15.5</points>
<intersection>-22 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>603,-22,650,-22</points>
<connection>
<GID>569</GID>
<name>IN_5</name></connection>
<intersection>603 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>556.5,-15.5,603,-15.5</points>
<connection>
<GID>641</GID>
<name>OUT</name></connection>
<intersection>603 0</intersection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>607,-60,607,-26.5</points>
<intersection>-60 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>607,-60,652,-60</points>
<connection>
<GID>454</GID>
<name>IN_5</name></connection>
<intersection>607 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>562,-26.5,607,-26.5</points>
<connection>
<GID>643</GID>
<name>OUT</name></connection>
<intersection>607 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>608.5,-37,608.5,-23</points>
<intersection>-37 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>608.5,-23,650,-23</points>
<connection>
<GID>569</GID>
<name>IN_4</name></connection>
<intersection>608.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>567,-37,608.5,-37</points>
<connection>
<GID>646</GID>
<name>OUT</name></connection>
<intersection>608.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>612,-61,612,-47</points>
<intersection>-61 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>612,-61,652,-61</points>
<connection>
<GID>454</GID>
<name>IN_4</name></connection>
<intersection>612 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>572.5,-47,612,-47</points>
<connection>
<GID>648</GID>
<name>OUT</name></connection>
<intersection>612 0</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>614,-57.5,614,-24</points>
<intersection>-57.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>614,-24,650,-24</points>
<connection>
<GID>569</GID>
<name>IN_3</name></connection>
<intersection>614 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>578,-57.5,614,-57.5</points>
<connection>
<GID>649</GID>
<name>OUT</name></connection>
<intersection>614 0</intersection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>617.5,-68,617.5,-62</points>
<intersection>-68 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>617.5,-62,652,-62</points>
<connection>
<GID>454</GID>
<name>IN_3</name></connection>
<intersection>617.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583.5,-68,617.5,-68</points>
<connection>
<GID>650</GID>
<name>OUT</name></connection>
<intersection>617.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>619,-78,619,-25</points>
<intersection>-78 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>619,-25,650,-25</points>
<connection>
<GID>569</GID>
<name>IN_2</name></connection>
<intersection>619 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588,-78,619,-78</points>
<connection>
<GID>572</GID>
<name>OUT</name></connection>
<intersection>619 0</intersection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>622.5,-88.5,622.5,-63</points>
<intersection>-88.5 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>622.5,-63,652,-63</points>
<connection>
<GID>454</GID>
<name>IN_2</name></connection>
<intersection>622.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>593.5,-88.5,622.5,-88.5</points>
<connection>
<GID>573</GID>
<name>OUT</name></connection>
<intersection>622.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493.5,-18.5,493.5,-12.5</points>
<intersection>-18.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,-18.5,493.5,-18.5</points>
<connection>
<GID>529</GID>
<name>OUT_5</name></connection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>493.5,-12.5,550.5,-12.5</points>
<connection>
<GID>641</GID>
<name>IN_3</name></connection>
<intersection>493.5 0</intersection>
<intersection>502.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>502.5,-23.5,502.5,-12.5</points>
<intersection>-23.5 4</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>502.5,-23.5,556,-23.5</points>
<connection>
<GID>643</GID>
<name>IN_3</name></connection>
<intersection>502.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495.5,-42.5,495.5,-14.5</points>
<intersection>-42.5 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>480,-42.5,495.5,-42.5</points>
<connection>
<GID>545</GID>
<name>OUT_5</name></connection>
<intersection>495.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>495.5,-14.5,550.5,-14.5</points>
<connection>
<GID>641</GID>
<name>IN_2</name></connection>
<intersection>495.5 0</intersection>
<intersection>504 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>504,-25.5,504,-14.5</points>
<intersection>-25.5 4</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>504,-25.5,556,-25.5</points>
<connection>
<GID>643</GID>
<name>IN_2</name></connection>
<intersection>504 3</intersection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>498,-67.5,498,-16.5</points>
<intersection>-67.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-67.5,498,-67.5</points>
<connection>
<GID>555</GID>
<name>OUT_5</name></connection>
<intersection>498 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>498,-16.5,550.5,-16.5</points>
<connection>
<GID>641</GID>
<name>IN_1</name></connection>
<intersection>498 0</intersection>
<intersection>506 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>506,-27.5,506,-16.5</points>
<intersection>-27.5 4</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>506,-27.5,556,-27.5</points>
<connection>
<GID>643</GID>
<name>IN_1</name></connection>
<intersection>506 3</intersection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>500.5,-92.5,500.5,-18.5</points>
<intersection>-92.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-92.5,500.5,-92.5</points>
<connection>
<GID>557</GID>
<name>OUT_5</name></connection>
<intersection>500.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>500.5,-18.5,550.5,-18.5</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>500.5 0</intersection>
<intersection>508.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>508.5,-29.5,508.5,-18.5</points>
<intersection>-29.5 4</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>508.5,-29.5,556,-29.5</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>508.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,-34,502,-19.5</points>
<intersection>-34 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,-19.5,502,-19.5</points>
<connection>
<GID>529</GID>
<name>OUT_4</name></connection>
<intersection>502 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>502,-34,561,-34</points>
<connection>
<GID>646</GID>
<name>IN_3</name></connection>
<intersection>502 0</intersection>
<intersection>509 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>509,-44,509,-34</points>
<intersection>-44 4</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>509,-44,566.5,-44</points>
<connection>
<GID>648</GID>
<name>IN_3</name></connection>
<intersection>509 3</intersection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502.5,-43.5,502.5,-36</points>
<intersection>-43.5 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>480,-43.5,502.5,-43.5</points>
<connection>
<GID>545</GID>
<name>OUT_4</name></connection>
<intersection>502.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>502.5,-36,561,-36</points>
<connection>
<GID>646</GID>
<name>IN_2</name></connection>
<intersection>502.5 0</intersection>
<intersection>511 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>511,-46,511,-36</points>
<intersection>-46 4</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>511,-46,566.5,-46</points>
<connection>
<GID>648</GID>
<name>IN_2</name></connection>
<intersection>511 3</intersection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>504.5,-68.5,504.5,-38</points>
<intersection>-68.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-68.5,504.5,-68.5</points>
<connection>
<GID>555</GID>
<name>OUT_4</name></connection>
<intersection>504.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>504.5,-38,561,-38</points>
<connection>
<GID>646</GID>
<name>IN_1</name></connection>
<intersection>504.5 0</intersection>
<intersection>513.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>513.5,-48,513.5,-38</points>
<intersection>-48 4</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>513.5,-48,566.5,-48</points>
<connection>
<GID>648</GID>
<name>IN_1</name></connection>
<intersection>513.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507,-93.5,507,-40</points>
<intersection>-93.5 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-93.5,507,-93.5</points>
<connection>
<GID>557</GID>
<name>OUT_4</name></connection>
<intersection>507 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>507,-40,561,-40</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>507 0</intersection>
<intersection>516 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>516,-50,516,-40</points>
<intersection>-50 4</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>516,-50,566.5,-50</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>516 3</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520,-54.5,520,-20.5</points>
<intersection>-54.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,-20.5,520,-20.5</points>
<connection>
<GID>529</GID>
<name>OUT_3</name></connection>
<intersection>520 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>520,-54.5,572,-54.5</points>
<connection>
<GID>649</GID>
<name>IN_3</name></connection>
<intersection>520 0</intersection>
<intersection>529 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>529,-65,529,-54.5</points>
<intersection>-65 4</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>529,-65,577.5,-65</points>
<connection>
<GID>650</GID>
<name>IN_3</name></connection>
<intersection>529 3</intersection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>521.5,-56.5,521.5,-44.5</points>
<intersection>-56.5 2</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>480,-44.5,521.5,-44.5</points>
<connection>
<GID>545</GID>
<name>OUT_3</name></connection>
<intersection>521.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>521.5,-56.5,572,-56.5</points>
<connection>
<GID>649</GID>
<name>IN_2</name></connection>
<intersection>521.5 0</intersection>
<intersection>531.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>531.5,-67,531.5,-56.5</points>
<intersection>-67 4</intersection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>531.5,-67,577.5,-67</points>
<connection>
<GID>650</GID>
<name>IN_2</name></connection>
<intersection>531.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>522.5,-69.5,522.5,-58.5</points>
<intersection>-69.5 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-69.5,522.5,-69.5</points>
<connection>
<GID>555</GID>
<name>OUT_3</name></connection>
<intersection>522.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>522.5,-58.5,572,-58.5</points>
<connection>
<GID>649</GID>
<name>IN_1</name></connection>
<intersection>522.5 0</intersection>
<intersection>534 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>534,-69,534,-58.5</points>
<intersection>-69 4</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>534,-69,577.5,-69</points>
<connection>
<GID>650</GID>
<name>IN_1</name></connection>
<intersection>534 3</intersection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524.5,-94.5,524.5,-60.5</points>
<intersection>-94.5 1</intersection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-94.5,524.5,-94.5</points>
<connection>
<GID>557</GID>
<name>OUT_3</name></connection>
<intersection>524.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>524.5,-60.5,572,-60.5</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>524.5 0</intersection>
<intersection>537 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>537,-71,537,-60.5</points>
<intersection>-71 4</intersection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>537,-71,577.5,-71</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>537 3</intersection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>559.5,-75,559.5,-21.5</points>
<intersection>-75 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,-21.5,559.5,-21.5</points>
<connection>
<GID>529</GID>
<name>OUT_2</name></connection>
<intersection>559.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>559.5,-75,582,-75</points>
<connection>
<GID>572</GID>
<name>IN_3</name></connection>
<intersection>559.5 0</intersection>
<intersection>563 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>563,-85.5,563,-75</points>
<intersection>-85.5 4</intersection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>563,-85.5,587.5,-85.5</points>
<connection>
<GID>573</GID>
<name>IN_3</name></connection>
<intersection>563 3</intersection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>557,-77,557,-45.5</points>
<intersection>-77 2</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>480,-45.5,557,-45.5</points>
<connection>
<GID>545</GID>
<name>OUT_2</name></connection>
<intersection>557 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>557,-77,582,-77</points>
<connection>
<GID>572</GID>
<name>IN_2</name></connection>
<intersection>557 0</intersection>
<intersection>565 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>565,-87.5,565,-77</points>
<intersection>-87.5 4</intersection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>565,-87.5,587.5,-87.5</points>
<connection>
<GID>573</GID>
<name>IN_2</name></connection>
<intersection>565 3</intersection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530.5,-79,530.5,-70.5</points>
<intersection>-79 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-70.5,530.5,-70.5</points>
<connection>
<GID>555</GID>
<name>OUT_2</name></connection>
<intersection>530.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>530.5,-79,582,-79</points>
<connection>
<GID>572</GID>
<name>IN_1</name></connection>
<intersection>530.5 0</intersection>
<intersection>567.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>567.5,-89.5,567.5,-79</points>
<intersection>-89.5 4</intersection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>567.5,-89.5,587.5,-89.5</points>
<connection>
<GID>573</GID>
<name>IN_1</name></connection>
<intersection>567.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530.5,-95.5,530.5,-81</points>
<intersection>-95.5 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-95.5,530.5,-95.5</points>
<connection>
<GID>557</GID>
<name>OUT_2</name></connection>
<intersection>530.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>530.5,-81,582,-81</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>530.5 0</intersection>
<intersection>569.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>569.5,-91.5,569.5,-81</points>
<intersection>-91.5 4</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>569.5,-91.5,587.5,-91.5</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>569.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>479.5,-16.5,479.5,26.5</points>
<intersection>-16.5 6</intersection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,26.5,525,26.5</points>
<connection>
<GID>645</GID>
<name>IN_3</name></connection>
<intersection>479.5 0</intersection>
<intersection>493 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>493,17,493,26.5</points>
<intersection>17 5</intersection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>493,17,531,17</points>
<connection>
<GID>664</GID>
<name>IN_3</name></connection>
<intersection>493 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>478.5,-16.5,479.5,-16.5</points>
<connection>
<GID>529</GID>
<name>OUT_7</name></connection>
<intersection>479.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>481,-40.5,481,24.5</points>
<intersection>-40.5 2</intersection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481,24.5,525,24.5</points>
<connection>
<GID>645</GID>
<name>IN_2</name></connection>
<intersection>481 0</intersection>
<intersection>491 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>480,-40.5,481,-40.5</points>
<connection>
<GID>545</GID>
<name>OUT_7</name></connection>
<intersection>481 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>491,15,491,24.5</points>
<intersection>15 4</intersection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>491,15,531,15</points>
<connection>
<GID>664</GID>
<name>IN_2</name></connection>
<intersection>491 3</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>483,-65.5,483,22.5</points>
<intersection>-65.5 2</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483,22.5,525,22.5</points>
<connection>
<GID>645</GID>
<name>IN_1</name></connection>
<intersection>483 0</intersection>
<intersection>489 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>479.5,-65.5,483,-65.5</points>
<connection>
<GID>555</GID>
<name>OUT_7</name></connection>
<intersection>483 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>489,13,489,22.5</points>
<intersection>13 4</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>489,13,531,13</points>
<connection>
<GID>664</GID>
<name>IN_1</name></connection>
<intersection>489 3</intersection></hsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616,-124,616,45.5</points>
<connection>
<GID>571</GID>
<name>SEL_0</name></connection>
<intersection>-83 11</intersection>
<intersection>-22.5 5</intersection>
<intersection>-4.5 3</intersection>
<intersection>45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>415.5,45.5,616,45.5</points>
<connection>
<GID>491</GID>
<name>OUT_0</name></connection>
<intersection>616 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>591.5,-4.5,616,-4.5</points>
<intersection>591.5 6</intersection>
<intersection>616 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>578,-22.5,616,-22.5</points>
<intersection>578 8</intersection>
<intersection>616 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>591.5,-4.5,591.5,19</points>
<intersection>-4.5 3</intersection>
<intersection>19 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>535,19,591.5,19</points>
<connection>
<GID>664</GID>
<name>SEL_0</name></connection>
<intersection>591.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>578,-22.5,578,0</points>
<intersection>-22.5 5</intersection>
<intersection>-21.5 12</intersection>
<intersection>0 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>548.5,0,578,0</points>
<intersection>548.5 10</intersection>
<intersection>578 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>548.5,-0.5,548.5,0</points>
<connection>
<GID>556</GID>
<name>SEL_0</name></connection>
<intersection>0 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>591.5,-83,616,-83</points>
<intersection>591.5 16</intersection>
<intersection>597 18</intersection>
<intersection>616 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>560,-21.5,581.5,-21.5</points>
<connection>
<GID>643</GID>
<name>SEL_0</name></connection>
<intersection>578 8</intersection>
<intersection>581.5 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>581.5,-63,581.5,-21.5</points>
<connection>
<GID>650</GID>
<name>SEL_0</name></connection>
<intersection>-40.5 15</intersection>
<intersection>-21.5 12</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>570.5,-40.5,581.5,-40.5</points>
<intersection>570.5 17</intersection>
<intersection>581.5 13</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>591.5,-83.5,591.5,-83</points>
<connection>
<GID>573</GID>
<name>SEL_0</name></connection>
<intersection>-83 11</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>570.5,-42,570.5,-40.5</points>
<connection>
<GID>648</GID>
<name>SEL_0</name></connection>
<intersection>-40.5 15</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>597,-94,597,-83</points>
<connection>
<GID>574</GID>
<name>SEL_0</name></connection>
<intersection>-83 11</intersection></vsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>588,4,588,49</points>
<intersection>4 5</intersection>
<intersection>20 9</intersection>
<intersection>49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>416,49,588,49</points>
<connection>
<GID>519</GID>
<name>OUT_0</name></connection>
<intersection>588 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>588,4,615,4</points>
<intersection>588 0</intersection>
<intersection>615 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>615,-124,615,4</points>
<connection>
<GID>571</GID>
<name>SEL_1</name></connection>
<intersection>-81.5 13</intersection>
<intersection>-25.5 8</intersection>
<intersection>4 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>574.5,-25.5,615,-25.5</points>
<intersection>574.5 10</intersection>
<intersection>580.5 18</intersection>
<intersection>615 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>534,20,588,20</points>
<intersection>534 15</intersection>
<intersection>588 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>574.5,-25.5,574.5,1.5</points>
<intersection>-25.5 8</intersection>
<intersection>-20 16</intersection>
<intersection>1.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>547.5,1.5,574.5,1.5</points>
<intersection>547.5 12</intersection>
<intersection>574.5 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>547.5,-0.5,547.5,1.5</points>
<connection>
<GID>556</GID>
<name>SEL_1</name></connection>
<intersection>1.5 11</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>590.5,-81.5,615,-81.5</points>
<intersection>590.5 21</intersection>
<intersection>596 14</intersection>
<intersection>615 6</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>596,-94,596,-81.5</points>
<connection>
<GID>574</GID>
<name>SEL_1</name></connection>
<intersection>-81.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>534,19,534,20</points>
<connection>
<GID>664</GID>
<name>SEL_1</name></connection>
<intersection>20 9</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>559,-20,574.5,-20</points>
<intersection>559 17</intersection>
<intersection>574.5 10</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>559,-21.5,559,-20</points>
<connection>
<GID>643</GID>
<name>SEL_1</name></connection>
<intersection>-20 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>580.5,-63,580.5,-25.5</points>
<connection>
<GID>650</GID>
<name>SEL_1</name></connection>
<intersection>-39.5 20</intersection>
<intersection>-25.5 8</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>569.5,-39.5,580.5,-39.5</points>
<intersection>569.5 22</intersection>
<intersection>580.5 18</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>590.5,-83.5,590.5,-81.5</points>
<connection>
<GID>573</GID>
<name>SEL_1</name></connection>
<intersection>-81.5 13</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>569.5,-42,569.5,-39.5</points>
<connection>
<GID>648</GID>
<name>SEL_1</name></connection>
<intersection>-39.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>528,28.5,528,35</points>
<connection>
<GID>645</GID>
<name>SEL_1</name></connection>
<intersection>35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>417,35,608,35</points>
<connection>
<GID>485</GID>
<name>OUT_0</name></connection>
<intersection>528 0</intersection>
<intersection>608 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>608,-114.5,608,35</points>
<connection>
<GID>570</GID>
<name>SEL_1</name></connection>
<intersection>-100.5 14</intersection>
<intersection>-13 8</intersection>
<intersection>35 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>580.5,-13,608,-13</points>
<intersection>580.5 9</intersection>
<intersection>608 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>580.5,-13,580.5,11.5</points>
<intersection>-13 8</intersection>
<intersection>11.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>541.5,11.5,585,11.5</points>
<intersection>541.5 16</intersection>
<intersection>580.5 9</intersection>
<intersection>585 17</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>601.5,-100.5,608,-100.5</points>
<intersection>601.5 15</intersection>
<intersection>608 6</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>601.5,-104,601.5,-100.5</points>
<connection>
<GID>575</GID>
<name>SEL_1</name></connection>
<intersection>-100.5 14</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>541.5,10.5,541.5,11.5</points>
<connection>
<GID>554</GID>
<name>SEL_1</name></connection>
<intersection>11.5 10</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>585,-73,585,11.5</points>
<connection>
<GID>572</GID>
<name>SEL_1</name></connection>
<intersection>-50.5 24</intersection>
<intersection>-29 22</intersection>
<intersection>-7.5 19</intersection>
<intersection>11.5 10</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>553.5,-7.5,585,-7.5</points>
<intersection>553.5 20</intersection>
<intersection>585 17</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>553.5,-10.5,553.5,-7.5</points>
<connection>
<GID>641</GID>
<name>SEL_1</name></connection>
<intersection>-7.5 19</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>564,-29,585,-29</points>
<intersection>564 25</intersection>
<intersection>585 17</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>575,-50.5,585,-50.5</points>
<intersection>575 26</intersection>
<intersection>585 17</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>564,-32,564,-29</points>
<connection>
<GID>646</GID>
<name>SEL_1</name></connection>
<intersection>-29 22</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>575,-52.5,575,-50.5</points>
<connection>
<GID>649</GID>
<name>SEL_1</name></connection>
<intersection>-50.5 24</intersection></vsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>393,-93.5,396.5,-93.5</points>
<connection>
<GID>651</GID>
<name>OUT_0</name></connection>
<intersection>396.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>396.5,-93.5,396.5,-87.5</points>
<intersection>-93.5 1</intersection>
<intersection>-87.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>396.5,-87.5,398.5,-87.5</points>
<connection>
<GID>662</GID>
<name>IN_1</name></connection>
<intersection>396.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397.5,-99.5,397.5,-88.5</points>
<intersection>-99.5 3</intersection>
<intersection>-88.5 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>387.5,-99.5,397.5,-99.5</points>
<intersection>387.5 6</intersection>
<intersection>397.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>397.5,-88.5,398.5,-88.5</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<intersection>397.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>387.5,-99.5,387.5,-99</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>-99.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>406,-14.5,473.5,-14.5</points>
<connection>
<GID>529</GID>
<name>load</name></connection>
<intersection>406 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>406,-85.5,406,-14.5</points>
<intersection>-85.5 7</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>404.5,-85.5,406,-85.5</points>
<connection>
<GID>662</GID>
<name>OUT_3</name></connection>
<intersection>406 3</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>148,-33,155.5,-33</points>
<connection>
<GID>470</GID>
<name>OUT_1</name></connection>
<connection>
<GID>495</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>148,-34,155.5,-34</points>
<connection>
<GID>470</GID>
<name>OUT_0</name></connection>
<connection>
<GID>495</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>146,-24.5,146,-22.5</points>
<intersection>-24.5 5</intersection>
<intersection>-22.5 11</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>143,-24.5,146,-24.5</points>
<intersection>143 7</intersection>
<intersection>146 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>143,-25,143,-24.5</points>
<connection>
<GID>470</GID>
<name>load</name></connection>
<intersection>-24.5 5</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>145.5,-22.5,146,-22.5</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<intersection>146 1</intersection></hsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,-35.5,226,-19.5</points>
<connection>
<GID>644</GID>
<name>DATA_OUT_10</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,-35.5,228.5,-35.5</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408,-86.5,408,-38.5</points>
<intersection>-86.5 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>404.5,-86.5,408,-86.5</points>
<connection>
<GID>662</GID>
<name>OUT_2</name></connection>
<intersection>408 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>408,-38.5,475,-38.5</points>
<connection>
<GID>545</GID>
<name>load</name></connection>
<intersection>408 0</intersection></hsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>202.5,59,203.5,59</points>
<connection>
<GID>479</GID>
<name>OUT_7</name></connection>
<connection>
<GID>480</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>202.5,58,203.5,58</points>
<connection>
<GID>479</GID>
<name>OUT_6</name></connection>
<connection>
<GID>480</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>202.5,57,203.5,57</points>
<connection>
<GID>479</GID>
<name>OUT_5</name></connection>
<connection>
<GID>480</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>202.5,56,203.5,56</points>
<connection>
<GID>479</GID>
<name>OUT_4</name></connection>
<connection>
<GID>480</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>202.5,55,203.5,55</points>
<connection>
<GID>479</GID>
<name>OUT_3</name></connection>
<connection>
<GID>480</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>202.5,54,203.5,54</points>
<connection>
<GID>479</GID>
<name>OUT_2</name></connection>
<connection>
<GID>480</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>202.5,53,203.5,53</points>
<connection>
<GID>479</GID>
<name>OUT_1</name></connection>
<connection>
<GID>480</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>202.5,52,203.5,52</points>
<connection>
<GID>479</GID>
<name>OUT_0</name></connection>
<connection>
<GID>480</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>199.5,46,199.5,50</points>
<connection>
<GID>481</GID>
<name>OUT_0</name></connection>
<connection>
<GID>479</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>26</ID>
<points>195,61,195,68.5</points>
<intersection>61 46</intersection>
<intersection>68.5 44</intersection></vsegment>
<hsegment>
<ID>44</ID>
<points>190.5,68.5,195,68.5</points>
<intersection>190.5 45</intersection>
<intersection>195 26</intersection></hsegment>
<vsegment>
<ID>45</ID>
<points>190.5,68.5,190.5,70.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>68.5 44</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>195,61,197.5,61</points>
<connection>
<GID>479</GID>
<name>load</name></connection>
<intersection>195 26</intersection></hsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-14.5,118.5,-8</points>
<intersection>-14.5 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,-14.5,121.5,-14.5</points>
<connection>
<GID>494</GID>
<name>ADDRESS_7</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-8,118.5,-8</points>
<intersection>92.5 3</intersection>
<intersection>118.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92.5,-8,92.5,-5</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<intersection>-8 2</intersection></vsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-15.5,117.5,-10.5</points>
<intersection>-15.5 1</intersection>
<intersection>-10.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-15.5,121.5,-15.5</points>
<connection>
<GID>494</GID>
<name>ADDRESS_6</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>92.5,-10.5,117.5,-10.5</points>
<intersection>92.5 4</intersection>
<intersection>117.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>92.5,-10.5,92.5,-9</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>-10.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-16.5,116.5,-12.5</points>
<intersection>-16.5 1</intersection>
<intersection>-12.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-16.5,121.5,-16.5</points>
<connection>
<GID>494</GID>
<name>ADDRESS_5</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>92.5,-12.5,116.5,-12.5</points>
<intersection>92.5 4</intersection>
<intersection>116.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>92.5,-12.5,92.5,-12</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>-12.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-17.5,115.5,-14.5</points>
<intersection>-17.5 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-17.5,121.5,-17.5</points>
<connection>
<GID>494</GID>
<name>ADDRESS_4</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-14.5,115.5,-14.5</points>
<intersection>92.5 3</intersection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92.5,-15,92.5,-14.5</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>-14.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-21.5,115.5,-18.5</points>
<intersection>-21.5 3</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-18.5,121.5,-18.5</points>
<connection>
<GID>494</GID>
<name>ADDRESS_3</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>92.5,-21.5,115.5,-21.5</points>
<intersection>92.5 4</intersection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>92.5,-21.5,92.5,-18.5</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>-21.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-23.5,116.5,-19.5</points>
<intersection>-23.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-19.5,121.5,-19.5</points>
<connection>
<GID>494</GID>
<name>ADDRESS_2</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-23.5,116.5,-23.5</points>
<intersection>92.5 3</intersection>
<intersection>116.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92.5,-23.5,92.5,-22</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>-23.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-25.5,117.5,-20.5</points>
<intersection>-25.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-20.5,121.5,-20.5</points>
<connection>
<GID>494</GID>
<name>ADDRESS_1</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-25.5,117.5,-25.5</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-27.5,118.5,-21.5</points>
<intersection>-27.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,-21.5,121.5,-21.5</points>
<connection>
<GID>494</GID>
<name>ADDRESS_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-27.5,118.5,-27.5</points>
<intersection>92.5 3</intersection>
<intersection>118.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92.5,-29,92.5,-27.5</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<intersection>-27.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,36.5,285.5,43.5</points>
<intersection>36.5 2</intersection>
<intersection>43.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>285.5,36.5,286.5,36.5</points>
<connection>
<GID>498</GID>
<name>IN_7</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281.5,43.5,285.5,43.5</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,35.5,284.5,40.5</points>
<intersection>35.5 1</intersection>
<intersection>40.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,35.5,286.5,35.5</points>
<connection>
<GID>498</GID>
<name>IN_6</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,40.5,284.5,40.5</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283.5,34.5,283.5,37.5</points>
<intersection>34.5 1</intersection>
<intersection>37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>283.5,34.5,286.5,34.5</points>
<connection>
<GID>498</GID>
<name>IN_5</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,37.5,283.5,37.5</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>282.5,33.5,282.5,34.5</points>
<intersection>33.5 8</intersection>
<intersection>34.5 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>282.5,33.5,286.5,33.5</points>
<connection>
<GID>498</GID>
<name>IN_4</name></connection>
<intersection>282.5 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>281.5,34.5,282.5,34.5</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<intersection>282.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,31.5,282.5,32.5</points>
<intersection>31.5 2</intersection>
<intersection>32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282.5,32.5,286.5,32.5</points>
<connection>
<GID>498</GID>
<name>IN_3</name></connection>
<intersection>282.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,31.5,282.5,31.5</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<intersection>282.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>281.5,28.5,283.5,28.5</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>283.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>283.5,28.5,283.5,31.5</points>
<intersection>28.5 1</intersection>
<intersection>31.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>283.5,31.5,286.5,31.5</points>
<connection>
<GID>498</GID>
<name>IN_2</name></connection>
<intersection>283.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,25.5,284.5,30.5</points>
<intersection>25.5 2</intersection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,30.5,286.5,30.5</points>
<connection>
<GID>498</GID>
<name>IN_1</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,25.5,284.5,25.5</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,22.5,285.5,29.5</points>
<intersection>22.5 2</intersection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>285.5,29.5,286.5,29.5</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,22.5,285.5,22.5</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,39.5,286,49</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>39.5 2</intersection>
<intersection>40.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>289.5,38.5,289.5,39.5</points>
<connection>
<GID>498</GID>
<name>load</name></connection>
<intersection>39.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>286,39.5,289.5,39.5</points>
<intersection>286 0</intersection>
<intersection>289.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>286,40.5,287.5,40.5</points>
<connection>
<GID>501</GID>
<name>OUT_0</name></connection>
<intersection>286 0</intersection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,33.5,295.5,58</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,33.5,316.5,33.5</points>
<connection>
<GID>498</GID>
<name>OUT_4</name></connection>
<connection>
<GID>510</GID>
<name>IN_4</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,34.5,296.5,58</points>
<connection>
<GID>520</GID>
<name>IN_1</name></connection>
<intersection>34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,34.5,316.5,34.5</points>
<connection>
<GID>498</GID>
<name>OUT_5</name></connection>
<connection>
<GID>510</GID>
<name>IN_5</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297.5,35.5,297.5,58</points>
<connection>
<GID>520</GID>
<name>IN_2</name></connection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,35.5,316.5,35.5</points>
<connection>
<GID>498</GID>
<name>OUT_6</name></connection>
<connection>
<GID>510</GID>
<name>IN_6</name></connection>
<intersection>297.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,36.5,298.5,58</points>
<connection>
<GID>520</GID>
<name>IN_3</name></connection>
<intersection>36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,36.5,316.5,36.5</points>
<connection>
<GID>498</GID>
<name>OUT_7</name></connection>
<connection>
<GID>510</GID>
<name>IN_7</name></connection>
<intersection>298.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315.5,32.5,315.5,58</points>
<connection>
<GID>521</GID>
<name>IN_3</name></connection>
<intersection>32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,32.5,316.5,32.5</points>
<connection>
<GID>498</GID>
<name>OUT_3</name></connection>
<connection>
<GID>510</GID>
<name>IN_3</name></connection>
<intersection>315.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,29.5,312.5,58</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,29.5,316.5,29.5</points>
<connection>
<GID>498</GID>
<name>OUT_0</name></connection>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>294.5,30.5,316.5,30.5</points>
<connection>
<GID>498</GID>
<name>OUT_1</name></connection>
<connection>
<GID>510</GID>
<name>IN_1</name></connection>
<intersection>313.5 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>313.5,30.5,313.5,58</points>
<connection>
<GID>521</GID>
<name>IN_1</name></connection>
<intersection>30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314.5,31.5,314.5,58</points>
<connection>
<GID>521</GID>
<name>IN_2</name></connection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,31.5,316.5,31.5</points>
<connection>
<GID>498</GID>
<name>OUT_2</name></connection>
<connection>
<GID>510</GID>
<name>IN_2</name></connection>
<intersection>314.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<hsegment>
<ID>13</ID>
<points>301.5,61,302.5,61</points>
<connection>
<GID>520</GID>
<name>carry_out</name></connection>
<connection>
<GID>521</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<hsegment>
<ID>13</ID>
<points>284.5,61,285.5,61</points>
<connection>
<GID>500</GID>
<name>OUT_0</name></connection>
<connection>
<GID>520</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>410,-87.5,410,-63.5</points>
<intersection>-87.5 1</intersection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>404.5,-87.5,410,-87.5</points>
<connection>
<GID>662</GID>
<name>OUT_1</name></connection>
<intersection>410 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>410,-63.5,474.5,-63.5</points>
<connection>
<GID>555</GID>
<name>load</name></connection>
<intersection>410 0</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,67,289,69</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>67 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>289,67,292,67</points>
<intersection>289 0</intersection>
<intersection>292 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>292,66,292,67</points>
<connection>
<GID>520</GID>
<name>OUT_0</name></connection>
<intersection>67 3</intersection></vsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,66,293,68</points>
<connection>
<GID>520</GID>
<name>OUT_1</name></connection>
<intersection>68 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>292,68,292,69</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<intersection>68 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>292,68,293,68</points>
<intersection>292 1</intersection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,66,294,68</points>
<connection>
<GID>520</GID>
<name>OUT_2</name></connection>
<intersection>68 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>294,68,295,68</points>
<intersection>294 0</intersection>
<intersection>295 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>295,68,295,69</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>68 3</intersection></vsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>295,67,298,67</points>
<intersection>295 4</intersection>
<intersection>298 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>295,66,295,67</points>
<connection>
<GID>520</GID>
<name>OUT_3</name></connection>
<intersection>67 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>298,67,298,69</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>67 3</intersection></vsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,68,309,69</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>68 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>310,66,310,68</points>
<connection>
<GID>521</GID>
<name>OUT_1</name></connection>
<intersection>68 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>309,68,310,68</points>
<intersection>309 0</intersection>
<intersection>310 1</intersection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,66,311,68</points>
<connection>
<GID>521</GID>
<name>OUT_2</name></connection>
<intersection>68 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>311,68,312,68</points>
<intersection>311 0</intersection>
<intersection>312 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>312,68,312,69</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>68 3</intersection></vsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>312,66,312,67</points>
<connection>
<GID>521</GID>
<name>OUT_3</name></connection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>312,67,315,67</points>
<intersection>312 1</intersection>
<intersection>315 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>315,67,315,69</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>67 2</intersection></vsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>309,66,309,67</points>
<connection>
<GID>521</GID>
<name>OUT_0</name></connection>
<intersection>67 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>306,67,309,67</points>
<intersection>306 3</intersection>
<intersection>309 1</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>306,67,306,69</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>67 2</intersection></vsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-47.5,130,-25</points>
<connection>
<GID>494</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>494</GID>
<name>DATA_IN_0</name></connection>
<intersection>-47.5 17</intersection>
<intersection>-34 28</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>121.5,-47.5,130,-47.5</points>
<connection>
<GID>524</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>130,-34,140,-34</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-46.5,129,-25</points>
<connection>
<GID>494</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>494</GID>
<name>DATA_IN_1</name></connection>
<intersection>-46.5 17</intersection>
<intersection>-33 46</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>121.5,-46.5,129,-46.5</points>
<connection>
<GID>524</GID>
<name>OUT_1</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>129,-33,140,-33</points>
<connection>
<GID>470</GID>
<name>IN_1</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-45.5,128,-25</points>
<connection>
<GID>494</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>494</GID>
<name>DATA_IN_2</name></connection>
<intersection>-45.5 10</intersection>
<intersection>-32 38</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>121.5,-45.5,128,-45.5</points>
<connection>
<GID>524</GID>
<name>OUT_2</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>128,-32,140,-32</points>
<connection>
<GID>470</GID>
<name>IN_2</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>127,-44.5,127,-25</points>
<connection>
<GID>494</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>494</GID>
<name>DATA_IN_3</name></connection>
<intersection>-44.5 20</intersection>
<intersection>-31 48</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>121.5,-44.5,127,-44.5</points>
<connection>
<GID>524</GID>
<name>OUT_3</name></connection>
<intersection>127 3</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>127,-31,140,-31</points>
<connection>
<GID>470</GID>
<name>IN_3</name></connection>
<intersection>127 3</intersection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-43.5,126,-25</points>
<connection>
<GID>494</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>494</GID>
<name>DATA_IN_4</name></connection>
<intersection>-43.5 17</intersection>
<intersection>-30 45</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>121.5,-43.5,126,-43.5</points>
<connection>
<GID>524</GID>
<name>OUT_4</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>126,-30,140,-30</points>
<connection>
<GID>470</GID>
<name>IN_4</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-42.5,125,-25</points>
<connection>
<GID>494</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>494</GID>
<name>DATA_IN_5</name></connection>
<intersection>-42.5 17</intersection>
<intersection>-29 31</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>121.5,-42.5,125,-42.5</points>
<connection>
<GID>524</GID>
<name>OUT_5</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>125,-29,140,-29</points>
<connection>
<GID>470</GID>
<name>IN_5</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-41.5,124,-25</points>
<connection>
<GID>494</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>494</GID>
<name>DATA_IN_6</name></connection>
<intersection>-41.5 46</intersection>
<intersection>-28 31</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>124,-28,140,-28</points>
<connection>
<GID>470</GID>
<name>IN_6</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>121.5,-41.5,124,-41.5</points>
<connection>
<GID>524</GID>
<name>OUT_6</name></connection>
<intersection>124 0</intersection></hsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-40.5,123,-25</points>
<connection>
<GID>494</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>494</GID>
<name>DATA_IN_7</name></connection>
<intersection>-40.5 10</intersection>
<intersection>-27 24</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>121.5,-40.5,123,-40.5</points>
<connection>
<GID>524</GID>
<name>OUT_7</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>123,-27,140,-27</points>
<connection>
<GID>470</GID>
<name>IN_7</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-26,132.5,-7.5</points>
<intersection>-26 3</intersection>
<intersection>-17.5 2</intersection>
<intersection>-7.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>131.5,-17.5,132.5,-17.5</points>
<connection>
<GID>494</GID>
<name>write_enable</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>119.5,-26,132.5,-26</points>
<intersection>119.5 4</intersection>
<intersection>132.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>119.5,-39,119.5,-26</points>
<connection>
<GID>524</GID>
<name>ENABLE_0</name></connection>
<intersection>-26 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>130.5,-7.5,132.5,-7.5</points>
<intersection>130.5 6</intersection>
<intersection>132.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>130.5,-7.5,130.5,-6</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<intersection>-7.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92,-34.5,116.5,-34.5</points>
<intersection>92 9</intersection>
<intersection>116.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,-40.5,116.5,-34.5</points>
<intersection>-40.5 6</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>116.5,-40.5,117.5,-40.5</points>
<connection>
<GID>524</GID>
<name>IN_7</name></connection>
<intersection>116.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>92,-34.5,92,-33.5</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>404.5,-88.5,474.5,-88.5</points>
<connection>
<GID>557</GID>
<name>load</name></connection>
<connection>
<GID>662</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>529,28.5,529,30.5</points>
<connection>
<GID>645</GID>
<name>SEL_0</name></connection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>417,30.5,609,30.5</points>
<connection>
<GID>482</GID>
<name>OUT_0</name></connection>
<intersection>529 0</intersection>
<intersection>609 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>609,-114.5,609,30.5</points>
<connection>
<GID>570</GID>
<name>SEL_0</name></connection>
<intersection>-101.5 13</intersection>
<intersection>-16 7</intersection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>584.5,-16,609,-16</points>
<intersection>584.5 8</intersection>
<intersection>609 5</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>584.5,-16,584.5,10.5</points>
<intersection>-16 7</intersection>
<intersection>10.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>542.5,10.5,586,10.5</points>
<connection>
<GID>554</GID>
<name>SEL_0</name></connection>
<intersection>584.5 8</intersection>
<intersection>586 15</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>602.5,-101.5,609,-101.5</points>
<intersection>602.5 14</intersection>
<intersection>609 5</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>602.5,-104,602.5,-101.5</points>
<connection>
<GID>575</GID>
<name>SEL_0</name></connection>
<intersection>-101.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>586,-73,586,10.5</points>
<connection>
<GID>572</GID>
<name>SEL_0</name></connection>
<intersection>-51.5 20</intersection>
<intersection>-30.5 16</intersection>
<intersection>-9 17</intersection>
<intersection>10.5 9</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>565,-30.5,586,-30.5</points>
<intersection>565 21</intersection>
<intersection>586 15</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>554.5,-9,586,-9</points>
<intersection>554.5 18</intersection>
<intersection>586 15</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>554.5,-10.5,554.5,-9</points>
<connection>
<GID>641</GID>
<name>SEL_0</name></connection>
<intersection>-9 17</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>576,-51.5,586,-51.5</points>
<intersection>576 22</intersection>
<intersection>586 15</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>565,-32,565,-30.5</points>
<connection>
<GID>646</GID>
<name>SEL_0</name></connection>
<intersection>-30.5 16</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>576,-52.5,576,-51.5</points>
<connection>
<GID>649</GID>
<name>SEL_0</name></connection>
<intersection>-51.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>596,-17.5,668.5,-17.5</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>596 8</intersection>
<intersection>650 11</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>596,-17.5,596,23.5</points>
<intersection>-17.5 1</intersection>
<intersection>23.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>531,23.5,596,23.5</points>
<connection>
<GID>645</GID>
<name>OUT</name></connection>
<intersection>596 8</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>650,-20,650,-17.5</points>
<connection>
<GID>569</GID>
<name>IN_7</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>390,-17.5,470.5,-17.5</points>
<connection>
<GID>529</GID>
<name>IN_6</name></connection>
<intersection>390 15</intersection>
<intersection>424 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>424,-41.5,424,-17.5</points>
<intersection>-41.5 6</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>424,-41.5,472,-41.5</points>
<connection>
<GID>545</GID>
<name>IN_6</name></connection>
<intersection>424 5</intersection>
<intersection>440 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>440,-66.5,440,-41.5</points>
<intersection>-66.5 9</intersection>
<intersection>-41.5 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>440,-66.5,471.5,-66.5</points>
<connection>
<GID>555</GID>
<name>IN_6</name></connection>
<intersection>440 8</intersection>
<intersection>456 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>456,-91.5,456,-66.5</points>
<intersection>-91.5 11</intersection>
<intersection>-66.5 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>456,-91.5,471.5,-91.5</points>
<connection>
<GID>557</GID>
<name>IN_6</name></connection>
<intersection>456 10</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>390,-23,390,-17.5</points>
<intersection>-23 16</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>380.5,-23,390,-23</points>
<intersection>380.5 20</intersection>
<intersection>390 15</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>380.5,-34,380.5,-23</points>
<intersection>-34 22</intersection>
<intersection>-23 16</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>379,-34,380.5,-34</points>
<connection>
<GID>450</GID>
<name>OUT_6</name></connection>
<intersection>380.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>115.5,-51.5,115.5,-46.5</points>
<intersection>-51.5 6</intersection>
<intersection>-46.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>115.5,-46.5,117.5,-46.5</points>
<connection>
<GID>524</GID>
<name>IN_1</name></connection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>92,-51.5,115.5,-51.5</points>
<intersection>92 9</intersection>
<intersection>115.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>92,-54,92,-51.5</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>-51.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-57.5,105,-47.5</points>
<intersection>-57.5 11</intersection>
<intersection>-47.5 12</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>92,-57.5,105,-57.5</points>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>105,-47.5,117.5,-47.5</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<hsegment>
<ID>20</ID>
<points>159.5,-27,175,-27</points>
<connection>
<GID>495</GID>
<name>OUT_7</name></connection>
<connection>
<GID>576</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>173,-29.5,173,-28</points>
<intersection>-29.5 18</intersection>
<intersection>-28 19</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>173,-29.5,174,-29.5</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>173 11</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>159.5,-28,173,-28</points>
<connection>
<GID>495</GID>
<name>OUT_6</name></connection>
<intersection>173 11</intersection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>172.5,-32,172.5,-29</points>
<intersection>-32 12</intersection>
<intersection>-29 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>172.5,-32,174,-32</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>172.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>159.5,-29,172.5,-29</points>
<connection>
<GID>495</GID>
<name>OUT_5</name></connection>
<intersection>172.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>171.5,-34.5,171.5,-30</points>
<intersection>-34.5 12</intersection>
<intersection>-30 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>171.5,-34.5,174,-34.5</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>171.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>159.5,-30,171.5,-30</points>
<connection>
<GID>495</GID>
<name>OUT_4</name></connection>
<intersection>171.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>171,-37.5,171,-31</points>
<intersection>-37.5 13</intersection>
<intersection>-31 14</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>171,-37.5,174,-37.5</points>
<connection>
<GID>620</GID>
<name>IN_0</name></connection>
<intersection>171 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>159.5,-31,171,-31</points>
<connection>
<GID>495</GID>
<name>OUT_3</name></connection>
<intersection>171 11</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>170.5,-40.5,170.5,-32</points>
<intersection>-40.5 12</intersection>
<intersection>-32 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>170.5,-40.5,174.5,-40.5</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>170.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>159.5,-32,170.5,-32</points>
<connection>
<GID>495</GID>
<name>OUT_2</name></connection>
<intersection>170.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>170,-43.5,170,-33</points>
<intersection>-43.5 12</intersection>
<intersection>-33 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>170,-43.5,174.5,-43.5</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>170 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>159.5,-33,170,-33</points>
<connection>
<GID>495</GID>
<name>OUT_1</name></connection>
<intersection>170 11</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<vsegment>
<ID>14</ID>
<points>169.5,-46.5,169.5,-34</points>
<intersection>-46.5 15</intersection>
<intersection>-34 16</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>169.5,-46.5,174.5,-46.5</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<intersection>169.5 14</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>159.5,-34,169.5,-34</points>
<connection>
<GID>495</GID>
<name>OUT_0</name></connection>
<intersection>169.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,60,127,62</points>
<connection>
<GID>530</GID>
<name>load</name></connection>
<connection>
<GID>532</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>129,47.5,129,49</points>
<connection>
<GID>534</GID>
<name>OUT_0</name></connection>
<connection>
<GID>530</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,39,116.5,51</points>
<intersection>39 2</intersection>
<intersection>51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,51,124,51</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,39,116.5,39</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,42.5,115,52</points>
<intersection>42.5 2</intersection>
<intersection>52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,52,124,52</points>
<connection>
<GID>530</GID>
<name>IN_1</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,42.5,115,42.5</points>
<connection>
<GID>543</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,47.5,113.5,53</points>
<intersection>47.5 2</intersection>
<intersection>53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,53,124,53</points>
<connection>
<GID>530</GID>
<name>IN_2</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,47.5,113.5,47.5</points>
<intersection>110 3</intersection>
<intersection>113.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,46,110,47.5</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>47.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,49.5,111.5,54</points>
<intersection>49.5 2</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,54,124,54</points>
<connection>
<GID>530</GID>
<name>IN_3</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,49.5,111.5,49.5</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,55,124,55</points>
<connection>
<GID>530</GID>
<name>IN_4</name></connection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,53,110,55</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>55 1</intersection></vsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,56,124,56</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<connection>
<GID>530</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,57,114,59.5</points>
<intersection>57 1</intersection>
<intersection>59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,57,124,57</points>
<connection>
<GID>530</GID>
<name>IN_6</name></connection>
<intersection>114 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,59.5,114,59.5</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,58,117.5,63</points>
<intersection>58 3</intersection>
<intersection>63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>110,63,117.5,63</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>117.5,58,124,58</points>
<connection>
<GID>530</GID>
<name>IN_7</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,58,132,64.5</points>
<connection>
<GID>530</GID>
<name>OUT_7</name></connection>
<intersection>64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,64.5,140.5,64.5</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,57,135.5,62</points>
<intersection>57 2</intersection>
<intersection>62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,62,140.5,62</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,57,135.5,57</points>
<connection>
<GID>530</GID>
<name>OUT_6</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,56,137.5,59.5</points>
<intersection>56 2</intersection>
<intersection>59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,59.5,140.5,59.5</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>137.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,56,137.5,56</points>
<connection>
<GID>530</GID>
<name>OUT_5</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,55,138.5,56.5</points>
<intersection>55 2</intersection>
<intersection>56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,56.5,140.5,56.5</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,55,138.5,55</points>
<connection>
<GID>530</GID>
<name>OUT_4</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>132,54,140.5,54</points>
<connection>
<GID>530</GID>
<name>OUT_3</name></connection>
<connection>
<GID>550</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,50.5,135,53</points>
<intersection>50.5 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,50.5,140.5,50.5</points>
<connection>
<GID>551</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,53,135,53</points>
<connection>
<GID>530</GID>
<name>OUT_2</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,47.5,134,52</points>
<intersection>47.5 1</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,47.5,140.5,47.5</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,52,134,52</points>
<connection>
<GID>530</GID>
<name>OUT_1</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,44.5,133,51</points>
<intersection>44.5 1</intersection>
<intersection>51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,44.5,140.5,44.5</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,51,133,51</points>
<connection>
<GID>530</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>392.5,-18.5,470.5,-18.5</points>
<connection>
<GID>529</GID>
<name>IN_5</name></connection>
<intersection>392.5 10</intersection>
<intersection>422 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>422,-42.5,422,-18.5</points>
<intersection>-42.5 9</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>422,-42.5,472,-42.5</points>
<connection>
<GID>545</GID>
<name>IN_5</name></connection>
<intersection>422 8</intersection>
<intersection>438 12</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>392.5,-28,392.5,-18.5</points>
<intersection>-28 11</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>381.5,-28,392.5,-28</points>
<intersection>381.5 19</intersection>
<intersection>392.5 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>438,-67.5,438,-42.5</points>
<intersection>-67.5 13</intersection>
<intersection>-42.5 9</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>438,-67.5,471.5,-67.5</points>
<connection>
<GID>555</GID>
<name>IN_5</name></connection>
<intersection>438 12</intersection>
<intersection>454 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>454,-92.5,454,-67.5</points>
<intersection>-92.5 15</intersection>
<intersection>-67.5 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>454,-92.5,471.5,-92.5</points>
<connection>
<GID>557</GID>
<name>IN_5</name></connection>
<intersection>454 14</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>381.5,-35,381.5,-28</points>
<intersection>-35 21</intersection>
<intersection>-28 11</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>379,-35,381.5,-35</points>
<connection>
<GID>450</GID>
<name>OUT_5</name></connection>
<intersection>381.5 19</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>394.5,-19.5,470.5,-19.5</points>
<connection>
<GID>529</GID>
<name>IN_4</name></connection>
<intersection>394.5 7</intersection>
<intersection>420 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>420,-43.5,420,-19.5</points>
<intersection>-43.5 6</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>420,-43.5,472,-43.5</points>
<connection>
<GID>545</GID>
<name>IN_4</name></connection>
<intersection>420 5</intersection>
<intersection>436 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>394.5,-30.5,394.5,-19.5</points>
<intersection>-30.5 8</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>382.5,-30.5,394.5,-30.5</points>
<intersection>382.5 16</intersection>
<intersection>394.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>436,-68.5,436,-43.5</points>
<intersection>-68.5 10</intersection>
<intersection>-43.5 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>436,-68.5,471.5,-68.5</points>
<connection>
<GID>555</GID>
<name>IN_4</name></connection>
<intersection>436 9</intersection>
<intersection>452 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>452,-93.5,452,-68.5</points>
<intersection>-93.5 12</intersection>
<intersection>-68.5 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>452,-93.5,471.5,-93.5</points>
<connection>
<GID>557</GID>
<name>IN_4</name></connection>
<intersection>452 11</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>382.5,-36,382.5,-30.5</points>
<intersection>-36 17</intersection>
<intersection>-30.5 8</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>379,-36,382.5,-36</points>
<connection>
<GID>450</GID>
<name>OUT_4</name></connection>
<intersection>382.5 16</intersection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>397,-20.5,470.5,-20.5</points>
<connection>
<GID>529</GID>
<name>IN_3</name></connection>
<intersection>397 7</intersection>
<intersection>418 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>418,-44.5,418,-20.5</points>
<intersection>-44.5 6</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>418,-44.5,472,-44.5</points>
<connection>
<GID>545</GID>
<name>IN_3</name></connection>
<intersection>418 5</intersection>
<intersection>434 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>397,-34,397,-20.5</points>
<intersection>-34 8</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>383.5,-34,397,-34</points>
<intersection>383.5 14</intersection>
<intersection>397 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>434,-69.5,434,-44.5</points>
<intersection>-69.5 10</intersection>
<intersection>-44.5 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>434,-69.5,471.5,-69.5</points>
<connection>
<GID>555</GID>
<name>IN_3</name></connection>
<intersection>434 9</intersection>
<intersection>450 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>450,-94.5,450,-69.5</points>
<intersection>-94.5 12</intersection>
<intersection>-69.5 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>450,-94.5,471.5,-94.5</points>
<connection>
<GID>557</GID>
<name>IN_3</name></connection>
<intersection>450 11</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>383.5,-37,383.5,-34</points>
<intersection>-37 15</intersection>
<intersection>-34 8</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>379,-37,383.5,-37</points>
<connection>
<GID>450</GID>
<name>OUT_3</name></connection>
<intersection>383.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>399,-21.5,470.5,-21.5</points>
<connection>
<GID>529</GID>
<name>IN_2</name></connection>
<intersection>399 7</intersection>
<intersection>416 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>416,-45.5,416,-21.5</points>
<intersection>-45.5 6</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>416,-45.5,472,-45.5</points>
<connection>
<GID>545</GID>
<name>IN_2</name></connection>
<intersection>416 5</intersection>
<intersection>432 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>399,-35,399,-21.5</points>
<intersection>-35 8</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>386.5,-35,399,-35</points>
<intersection>386.5 14</intersection>
<intersection>399 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>432,-70.5,432,-45.5</points>
<intersection>-70.5 10</intersection>
<intersection>-45.5 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>432,-70.5,471.5,-70.5</points>
<connection>
<GID>555</GID>
<name>IN_2</name></connection>
<intersection>432 9</intersection>
<intersection>448 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>448,-95.5,448,-70.5</points>
<intersection>-95.5 12</intersection>
<intersection>-70.5 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>448,-95.5,471.5,-95.5</points>
<connection>
<GID>557</GID>
<name>IN_2</name></connection>
<intersection>448 11</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>386.5,-38,386.5,-35</points>
<intersection>-38 17</intersection>
<intersection>-35 8</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>379,-38,386.5,-38</points>
<connection>
<GID>450</GID>
<name>OUT_2</name></connection>
<intersection>386.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>401,-22.5,470.5,-22.5</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>401 7</intersection>
<intersection>414 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>414,-46.5,414,-22.5</points>
<intersection>-46.5 6</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>414,-46.5,472,-46.5</points>
<connection>
<GID>545</GID>
<name>IN_1</name></connection>
<intersection>414 5</intersection>
<intersection>430 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>401,-39,401,-22.5</points>
<intersection>-39 8</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>379,-39,401,-39</points>
<connection>
<GID>450</GID>
<name>OUT_1</name></connection>
<intersection>401 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>430,-71.5,430,-46.5</points>
<intersection>-71.5 10</intersection>
<intersection>-46.5 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>430,-71.5,471.5,-71.5</points>
<connection>
<GID>555</GID>
<name>IN_1</name></connection>
<intersection>430 9</intersection>
<intersection>446 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>446,-96.5,446,-71.5</points>
<intersection>-96.5 12</intersection>
<intersection>-71.5 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>446,-96.5,471.5,-96.5</points>
<connection>
<GID>557</GID>
<name>IN_1</name></connection>
<intersection>446 11</intersection></hsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412,-23.5,470.5,-23.5</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>412 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>412,-47.5,412,-23.5</points>
<intersection>-47.5 6</intersection>
<intersection>-45.5 16</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>412,-47.5,472,-47.5</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<intersection>412 5</intersection>
<intersection>428 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>428,-72.5,428,-47.5</points>
<intersection>-72.5 10</intersection>
<intersection>-47.5 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>428,-72.5,471.5,-72.5</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>428 9</intersection>
<intersection>444 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>444,-97.5,444,-72.5</points>
<intersection>-97.5 12</intersection>
<intersection>-72.5 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>444,-97.5,471.5,-97.5</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>444 11</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>391,-45.5,412,-45.5</points>
<intersection>391 17</intersection>
<intersection>412 5</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>391,-45.5,391,-40</points>
<intersection>-45.5 16</intersection>
<intersection>-40 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>379,-40,391,-40</points>
<connection>
<GID>450</GID>
<name>OUT_0</name></connection>
<intersection>391 17</intersection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,59,192.5,66</points>
<intersection>59 2</intersection>
<intersection>66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,66,192.5,66</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>192.5,59,194.5,59</points>
<connection>
<GID>479</GID>
<name>IN_7</name></connection>
<intersection>192.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,58,190.5,62.5</points>
<intersection>58 1</intersection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190.5,58,194.5,58</points>
<connection>
<GID>479</GID>
<name>IN_6</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189.5,62.5,190.5,62.5</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,57,194.5,57</points>
<connection>
<GID>479</GID>
<name>IN_5</name></connection>
<intersection>189 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>189,57,189,59</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>57 1</intersection></vsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,56,194.5,56</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<connection>
<GID>479</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,52.5,190.5,55</points>
<intersection>52.5 2</intersection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190.5,55,194.5,55</points>
<connection>
<GID>479</GID>
<name>IN_3</name></connection>
<intersection>190.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,52.5,190.5,52.5</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,49,191.5,54</points>
<intersection>49 2</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,54,194.5,54</points>
<connection>
<GID>479</GID>
<name>IN_2</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,49,191.5,49</points>
<connection>
<GID>566</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,45.5,192.5,53</points>
<intersection>45.5 2</intersection>
<intersection>53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192.5,53,194.5,53</points>
<connection>
<GID>479</GID>
<name>IN_1</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,45.5,192.5,45.5</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,42,191.5,52</points>
<intersection>42 7</intersection>
<intersection>52 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>189,42,191.5,42</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>191.5,52,194.5,52</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>379,-16.5,470.5,-16.5</points>
<connection>
<GID>529</GID>
<name>IN_7</name></connection>
<intersection>379 20</intersection>
<intersection>426 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>426,-40.5,426,-16.5</points>
<intersection>-40.5 4</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>426,-40.5,472,-40.5</points>
<connection>
<GID>545</GID>
<name>IN_7</name></connection>
<intersection>426 3</intersection>
<intersection>442 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>442,-65.5,442,-40.5</points>
<intersection>-65.5 6</intersection>
<intersection>-40.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>442,-65.5,471.5,-65.5</points>
<connection>
<GID>555</GID>
<name>IN_7</name></connection>
<intersection>442 5</intersection>
<intersection>458 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>458,-90.5,458,-65.5</points>
<intersection>-90.5 8</intersection>
<intersection>-65.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>458,-90.5,471.5,-90.5</points>
<connection>
<GID>557</GID>
<name>IN_7</name></connection>
<intersection>458 7</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>379,-33,379,-16.5</points>
<connection>
<GID>450</GID>
<name>OUT_7</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>598,-55.5,598,14</points>
<intersection>-55.5 1</intersection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>598,-55.5,670.5,-55.5</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>598 0</intersection>
<intersection>652 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>537,14,598,14</points>
<connection>
<GID>664</GID>
<name>OUT</name></connection>
<intersection>598 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>652,-58,652,-55.5</points>
<connection>
<GID>454</GID>
<name>IN_7</name></connection>
<intersection>-55.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,19.5,122.5,49</points>
<intersection>19.5 3</intersection>
<intersection>49 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>122.5,49,127,49</points>
<connection>
<GID>530</GID>
<name>clock</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>122.5,19.5,289.5,19.5</points>
<intersection>122.5 0</intersection>
<intersection>168 6</intersection>
<intersection>177 4</intersection>
<intersection>197.5 8</intersection>
<intersection>289.5 7</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>177,-16.5,177,19.5</points>
<intersection>-16.5 5</intersection>
<intersection>19.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>131.5,-16.5,177,-16.5</points>
<connection>
<GID>494</GID>
<name>write_clock</name></connection>
<intersection>152.5 9</intersection>
<intersection>177 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>168,19.5,168,24.5</points>
<connection>
<GID>624</GID>
<name>CLK</name></connection>
<intersection>19.5 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>289.5,-77.5,289.5,27.5</points>
<connection>
<GID>498</GID>
<name>clock</name></connection>
<intersection>-77.5 15</intersection>
<intersection>-52.5 14</intersection>
<intersection>-27.5 17</intersection>
<intersection>-4 19</intersection>
<intersection>19.5 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>197.5,19.5,197.5,50</points>
<connection>
<GID>479</GID>
<name>clock</name></connection>
<intersection>19.5 3</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>152.5,-36,152.5,-16.5</points>
<intersection>-36 10</intersection>
<intersection>-16.5 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>143,-36,152.5,-36</points>
<connection>
<GID>470</GID>
<name>clock</name></connection>
<intersection>152.5 9</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>289.5,-52.5,474.5,-52.5</points>
<intersection>289.5 7</intersection>
<intersection>474.5 24</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>289.5,-77.5,474.5,-77.5</points>
<intersection>289.5 7</intersection>
<intersection>474.5 24</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>289.5,-27.5,475,-27.5</points>
<intersection>289.5 7</intersection>
<intersection>475 23</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>289.5,-4,473.5,-4</points>
<intersection>289.5 7</intersection>
<intersection>473.5 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>473.5,-25.5,473.5,-4</points>
<connection>
<GID>529</GID>
<name>clock</name></connection>
<intersection>-4 19</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>475,-49.5,475,-27.5</points>
<connection>
<GID>545</GID>
<name>clock</name></connection>
<intersection>-27.5 17</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>474.5,-99.5,474.5,-52.5</points>
<connection>
<GID>555</GID>
<name>clock</name></connection>
<connection>
<GID>557</GID>
<name>clock</name></connection>
<intersection>-77.5 15</intersection>
<intersection>-52.5 14</intersection></vsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-41.5,104.5,-37.5</points>
<intersection>-41.5 1</intersection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-41.5,117.5,-41.5</points>
<connection>
<GID>524</GID>
<name>IN_6</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-37.5,104.5,-37.5</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-42.5,105,-40.5</points>
<intersection>-42.5 1</intersection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-42.5,117.5,-42.5</points>
<connection>
<GID>524</GID>
<name>IN_5</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,-40.5,105,-40.5</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92,-43.5,117.5,-43.5</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<connection>
<GID>524</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>480,8.5,538.5,8.5</points>
<connection>
<GID>554</GID>
<name>IN_3</name></connection>
<intersection>480 8</intersection>
<intersection>500 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>500,-2.5,500,8.5</points>
<intersection>-2.5 4</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>500,-2.5,544.5,-2.5</points>
<connection>
<GID>556</GID>
<name>IN_3</name></connection>
<intersection>500 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>480,-17.5,480,8.5</points>
<intersection>-17.5 9</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>478.5,-17.5,480,-17.5</points>
<connection>
<GID>529</GID>
<name>OUT_6</name></connection>
<intersection>480 8</intersection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-45.5,117.5,-45.5</points>
<connection>
<GID>524</GID>
<name>IN_2</name></connection>
<intersection>98 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>98,-50.5,98,-45.5</points>
<intersection>-50.5 6</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>92,-50.5,98,-50.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>98 3</intersection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92,-47,117.5,-47</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>117.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>117.5,-47,117.5,-44.5</points>
<connection>
<GID>524</GID>
<name>IN_3</name></connection>
<intersection>-47 1</intersection></vsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322.5,22.5,322.5,29.5</points>
<intersection>22.5 1</intersection>
<intersection>29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322.5,22.5,335,22.5</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>322.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>320.5,29.5,322.5,29.5</points>
<connection>
<GID>510</GID>
<name>OUT_0</name></connection>
<intersection>322.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323.5,27.5,323.5,30.5</points>
<intersection>27.5 1</intersection>
<intersection>30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323.5,27.5,335,27.5</points>
<intersection>323.5 0</intersection>
<intersection>335 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>320.5,30.5,323.5,30.5</points>
<connection>
<GID>510</GID>
<name>OUT_1</name></connection>
<intersection>323.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>335,25.5,335,27.5</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322,38,322,49</points>
<intersection>38 2</intersection>
<intersection>49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,49,328.5,49</points>
<intersection>322 0</intersection>
<intersection>328.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>318.5,38,322,38</points>
<connection>
<GID>510</GID>
<name>ENABLE_0</name></connection>
<intersection>322 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>328.5,49,328.5,53</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>49 1</intersection></vsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325,28.5,325,31.5</points>
<intersection>28.5 2</intersection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,31.5,325,31.5</points>
<connection>
<GID>510</GID>
<name>OUT_2</name></connection>
<intersection>325 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>325,28.5,335,28.5</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>325 0</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,31.5,327.5,32.5</points>
<intersection>31.5 1</intersection>
<intersection>32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327.5,31.5,334.5,31.5</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>327.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>320.5,32.5,327.5,32.5</points>
<connection>
<GID>510</GID>
<name>OUT_3</name></connection>
<intersection>327.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,33.5,329.5,34.5</points>
<intersection>33.5 1</intersection>
<intersection>34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,33.5,329.5,33.5</points>
<connection>
<GID>510</GID>
<name>OUT_4</name></connection>
<intersection>329.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>329.5,34.5,334.5,34.5</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>329.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329,34.5,329,37</points>
<intersection>34.5 2</intersection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>329,37,334.5,37</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>329 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>320.5,34.5,329,34.5</points>
<connection>
<GID>510</GID>
<name>OUT_5</name></connection>
<intersection>329 0</intersection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,35.5,327.5,39.5</points>
<intersection>35.5 1</intersection>
<intersection>39.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,35.5,327.5,35.5</points>
<connection>
<GID>510</GID>
<name>OUT_6</name></connection>
<intersection>327.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>327.5,39.5,334.5,39.5</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>327.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326,36.5,326,42</points>
<intersection>36.5 2</intersection>
<intersection>42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>326,42,335.5,42</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>320.5,36.5,326,36.5</points>
<connection>
<GID>510</GID>
<name>OUT_7</name></connection>
<intersection>326 0</intersection></hsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>487,6.5,538.5,6.5</points>
<connection>
<GID>554</GID>
<name>IN_2</name></connection>
<intersection>487 5</intersection>
<intersection>498 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>498,-4.5,498,6.5</points>
<intersection>-4.5 4</intersection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>498,-4.5,544.5,-4.5</points>
<connection>
<GID>556</GID>
<name>IN_2</name></connection>
<intersection>498 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>487,-41.5,487,6.5</points>
<intersection>-41.5 6</intersection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>480,-41.5,487,-41.5</points>
<connection>
<GID>545</GID>
<name>OUT_6</name></connection>
<intersection>487 5</intersection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>489,-66.5,489,4.5</points>
<intersection>-66.5 1</intersection>
<intersection>4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-66.5,489,-66.5</points>
<connection>
<GID>555</GID>
<name>OUT_6</name></connection>
<intersection>489 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>489,4.5,538.5,4.5</points>
<connection>
<GID>554</GID>
<name>IN_1</name></connection>
<intersection>489 0</intersection>
<intersection>496 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>496,-6.5,496,4.5</points>
<intersection>-6.5 4</intersection>
<intersection>4.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>496,-6.5,544.5,-6.5</points>
<connection>
<GID>556</GID>
<name>IN_1</name></connection>
<intersection>496 3</intersection></hsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,-11,213.5,57</points>
<intersection>-11 1</intersection>
<intersection>57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-11,219.5,-11</points>
<connection>
<GID>644</GID>
<name>ADDRESS_3</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207.5,57,213.5,57</points>
<connection>
<GID>480</GID>
<name>OUT_5</name></connection>
<intersection>213.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>485,-90.5,485,20.5</points>
<intersection>-90.5 1</intersection>
<intersection>20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-90.5,485,-90.5</points>
<connection>
<GID>557</GID>
<name>OUT_7</name></connection>
<intersection>485 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>485,20.5,525,20.5</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>485 0</intersection>
<intersection>487 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>487,11,487,20.5</points>
<intersection>11 4</intersection>
<intersection>20.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>487,11,531,11</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<intersection>487 3</intersection></hsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221,-54,221,-19.5</points>
<connection>
<GID>644</GID>
<name>DATA_OUT_15</name></connection>
<intersection>-54 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>221,-54,221.5,-54</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>221 0</intersection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-50.5,222,-19.5</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<connection>
<GID>644</GID>
<name>DATA_OUT_14</name></connection></vsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-42,224,-19.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<connection>
<GID>644</GID>
<name>DATA_OUT_12</name></connection></vsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,-46.5,223,-19.5</points>
<connection>
<GID>644</GID>
<name>DATA_OUT_13</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223,-46.5,223.5,-46.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>223 0</intersection></hsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,-91.5,491.5,2.5</points>
<intersection>-91.5 1</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-91.5,491.5,-91.5</points>
<connection>
<GID>557</GID>
<name>OUT_6</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>491.5,2.5,538.5,2.5</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>491.5 0</intersection>
<intersection>494 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>494,-8.5,494,2.5</points>
<intersection>-8.5 4</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>494,-8.5,544.5,-8.5</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>494 3</intersection></hsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>544.5,5.5,637,5.5</points>
<connection>
<GID>554</GID>
<name>OUT</name></connection>
<intersection>637 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>637,-21,637,5.5</points>
<intersection>-21 5</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>637,-21,650,-21</points>
<connection>
<GID>569</GID>
<name>IN_6</name></connection>
<intersection>637 4</intersection></hsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596.5,-53.5,596.5,-5.5</points>
<intersection>-53.5 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>596.5,-53.5,667.5,-53.5</points>
<intersection>596.5 0</intersection>
<intersection>650.5 4</intersection>
<intersection>667.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>550.5,-5.5,596.5,-5.5</points>
<connection>
<GID>556</GID>
<name>OUT</name></connection>
<intersection>596.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>667.5,-58.5,667.5,-53.5</points>
<intersection>-58.5 6</intersection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>650.5,-59,650.5,-53.5</points>
<intersection>-59 5</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>650.5,-59,652,-59</points>
<connection>
<GID>454</GID>
<name>IN_6</name></connection>
<intersection>650.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>667.5,-58.5,670.5,-58.5</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>667.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>479.5,-132,612,-132</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>479.5 6</intersection>
<intersection>603.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>603.5,-132,603.5,-122.5</points>
<intersection>-132 1</intersection>
<intersection>-122.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>603.5,-122.5,605,-122.5</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<intersection>603.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>479.5,-132,479.5,-97.5</points>
<connection>
<GID>557</GID>
<name>OUT_0</name></connection>
<intersection>-132 1</intersection></vsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>525,-130,525,-72.5</points>
<intersection>-130 1</intersection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,-130,612,-130</points>
<connection>
<GID>571</GID>
<name>IN_1</name></connection>
<intersection>525 0</intersection>
<intersection>601.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>479.5,-72.5,525,-72.5</points>
<connection>
<GID>555</GID>
<name>OUT_0</name></connection>
<intersection>525 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>601.5,-130,601.5,-120.5</points>
<intersection>-130 1</intersection>
<intersection>-120.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>601.5,-120.5,605,-120.5</points>
<connection>
<GID>570</GID>
<name>IN_1</name></connection>
<intersection>601.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-10,214.5,58</points>
<intersection>-10 1</intersection>
<intersection>58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214.5,-10,219.5,-10</points>
<connection>
<GID>644</GID>
<name>ADDRESS_4</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207.5,58,214.5,58</points>
<connection>
<GID>480</GID>
<name>OUT_6</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,-9,215.5,59</points>
<intersection>-9 1</intersection>
<intersection>59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-9,219.5,-9</points>
<connection>
<GID>644</GID>
<name>ADDRESS_5</name></connection>
<intersection>215.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207.5,59,215.5,59</points>
<connection>
<GID>480</GID>
<name>OUT_7</name></connection>
<intersection>215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212.5,60.5,212.5,66</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>205.5,60.5,212.5,60.5</points>
<connection>
<GID>480</GID>
<name>ENABLE_0</name></connection>
<intersection>212.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-33,227,-19.5</points>
<connection>
<GID>644</GID>
<name>DATA_OUT_9</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,-33,228.5,-33</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,32,218,47.5</points>
<intersection>32 1</intersection>
<intersection>47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,32,226.5,32</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207.5,47.5,218,47.5</points>
<intersection>207.5 3</intersection>
<intersection>218 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>207.5,47.5,207.5,52</points>
<connection>
<GID>480</GID>
<name>OUT_0</name></connection>
<intersection>47.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220.5,35,220.5,48.5</points>
<intersection>35 1</intersection>
<intersection>48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220.5,35,226.5,35</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<intersection>220.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>208.5,48.5,220.5,48.5</points>
<intersection>208.5 3</intersection>
<intersection>220.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>208.5,48.5,208.5,53</points>
<intersection>48.5 2</intersection>
<intersection>53 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>207.5,53,208.5,53</points>
<connection>
<GID>480</GID>
<name>OUT_1</name></connection>
<intersection>208.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221.5,38,221.5,50</points>
<intersection>38 2</intersection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210,50,221.5,50</points>
<intersection>210 3</intersection>
<intersection>221.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>221.5,38,226.5,38</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>221.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>210,50,210,54</points>
<intersection>50 1</intersection>
<intersection>54 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>207.5,54,210,54</points>
<connection>
<GID>480</GID>
<name>OUT_2</name></connection>
<intersection>210 3</intersection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207.5,55,212.5,55</points>
<connection>
<GID>480</GID>
<name>OUT_3</name></connection>
<intersection>212.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>212.5,51,212.5,55</points>
<intersection>51 4</intersection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>212.5,51,223,51</points>
<intersection>212.5 3</intersection>
<intersection>223 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>223,41,223,51</points>
<intersection>41 6</intersection>
<intersection>51 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>223,41,226,41</points>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<intersection>223 5</intersection></hsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224.5,44,224.5,53.5</points>
<intersection>44 2</intersection>
<intersection>46.5 3</intersection>
<intersection>49 4</intersection>
<intersection>51.5 5</intersection>
<intersection>53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223.5,53.5,224.5,53.5</points>
<connection>
<GID>581</GID>
<name>OUT_0</name></connection>
<intersection>224.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>224.5,44,226,44</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>224.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>224.5,46.5,226,46.5</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>224.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>224.5,49,226,49</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>224.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>224.5,51.5,227,51.5</points>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<intersection>224.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-25.5,236,-19.5</points>
<connection>
<GID>644</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-25.5,236,-25.5</points>
<intersection>218 2</intersection>
<intersection>236 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>218,-25.5,218,-14</points>
<intersection>-25.5 1</intersection>
<intersection>-14 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>218,-14,219.5,-14</points>
<connection>
<GID>644</GID>
<name>ADDRESS_0</name></connection>
<intersection>218 2</intersection></hsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,-25,235,-19.5</points>
<connection>
<GID>644</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216.5,-25,235,-25</points>
<intersection>216.5 2</intersection>
<intersection>235 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>216.5,-25,216.5,-13</points>
<intersection>-25 1</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216.5,-13,219.5,-13</points>
<connection>
<GID>644</GID>
<name>ADDRESS_1</name></connection>
<intersection>216.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215,-23,215,-12</points>
<intersection>-23 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215,-12,219.5,-12</points>
<connection>
<GID>644</GID>
<name>ADDRESS_2</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>215,-23,234,-23</points>
<intersection>215 0</intersection>
<intersection>234 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>234,-23,234,-19.5</points>
<connection>
<GID>644</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-23 2</intersection></vsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369.5,-85.5,369.5,-9.5</points>
<intersection>-85.5 2</intersection>
<intersection>-31.5 3</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>369.5,-9.5,371.5,-9.5</points>
<connection>
<GID>590</GID>
<name>IN_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>369.5,-85.5,398.5,-85.5</points>
<connection>
<GID>662</GID>
<name>ENABLE</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>369.5,-31.5,377,-31.5</points>
<connection>
<GID>450</GID>
<name>ENABLE_0</name></connection>
<intersection>369.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-30,228,-19.5</points>
<connection>
<GID>644</GID>
<name>DATA_OUT_8</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228,-30,231,-30</points>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>309.5,-142.5,309.5,-142.5</points>
<connection>
<GID>616</GID>
<name>carry_out</name></connection>
<connection>
<GID>617</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-155.5,290,-127.5</points>
<intersection>-155.5 1</intersection>
<intersection>-127.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-155.5,306.5,-155.5</points>
<connection>
<GID>617</GID>
<name>IN_3</name></connection>
<intersection>290 0</intersection>
<intersection>306.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-127.5,290,-127.5</points>
<connection>
<GID>618</GID>
<name>OUT_3</name></connection>
<intersection>290 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>306.5,-160,306.5,-155.5</points>
<intersection>-160 4</intersection>
<intersection>-155.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>306.5,-160,307,-160</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<intersection>306.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-154.5,289,-129.5</points>
<intersection>-154.5 1</intersection>
<intersection>-129.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,-154.5,306.5,-154.5</points>
<connection>
<GID>617</GID>
<name>IN_2</name></connection>
<intersection>289 0</intersection>
<intersection>306.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-129.5,289,-129.5</points>
<connection>
<GID>618</GID>
<name>OUT_2</name></connection>
<intersection>289 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>306.5,-165.5,306.5,-154.5</points>
<intersection>-165.5 4</intersection>
<intersection>-154.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>306.5,-165.5,307,-165.5</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<intersection>306.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-153.5,288,-131.5</points>
<intersection>-153.5 1</intersection>
<intersection>-131.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288,-153.5,306.5,-153.5</points>
<connection>
<GID>617</GID>
<name>IN_1</name></connection>
<intersection>288 0</intersection>
<intersection>306 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-131.5,288,-131.5</points>
<connection>
<GID>618</GID>
<name>OUT_1</name></connection>
<intersection>288 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>306,-171,306,-153.5</points>
<intersection>-171 4</intersection>
<intersection>-153.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>306,-171,307,-171</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>306 3</intersection></hsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-152.5,287,-133.5</points>
<intersection>-152.5 1</intersection>
<intersection>-133.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-152.5,306.5,-152.5</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>287 0</intersection>
<intersection>306 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-133.5,287,-133.5</points>
<connection>
<GID>618</GID>
<name>OUT_0</name></connection>
<intersection>287 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>306,-176.5,306,-152.5</points>
<intersection>-176.5 4</intersection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>306,-176.5,307,-176.5</points>
<connection>
<GID>598</GID>
<name>IN_0</name></connection>
<intersection>306 3</intersection></hsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-156,290.5,-148.5</points>
<intersection>-156 2</intersection>
<intersection>-148.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,-148.5,306.5,-148.5</points>
<connection>
<GID>617</GID>
<name>IN_B_3</name></connection>
<intersection>290.5 0</intersection>
<intersection>306.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-156,290.5,-156</points>
<connection>
<GID>593</GID>
<name>OUT_3</name></connection>
<intersection>290.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>306.5,-162,306.5,-148.5</points>
<intersection>-162 4</intersection>
<intersection>-148.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>306.5,-162,307,-162</points>
<connection>
<GID>595</GID>
<name>IN_1</name></connection>
<intersection>306.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289.5,-167.5,289.5,-147.5</points>
<intersection>-167.5 3</intersection>
<intersection>-158 2</intersection>
<intersection>-147.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289.5,-147.5,306.5,-147.5</points>
<connection>
<GID>617</GID>
<name>IN_B_2</name></connection>
<intersection>289.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-158,289.5,-158</points>
<connection>
<GID>593</GID>
<name>OUT_2</name></connection>
<intersection>289.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>289.5,-167.5,307,-167.5</points>
<connection>
<GID>596</GID>
<name>IN_1</name></connection>
<intersection>289.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-173,288.5,-146.5</points>
<intersection>-173 3</intersection>
<intersection>-160 2</intersection>
<intersection>-146.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288.5,-146.5,306.5,-146.5</points>
<connection>
<GID>617</GID>
<name>IN_B_1</name></connection>
<intersection>288.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-160,288.5,-160</points>
<connection>
<GID>593</GID>
<name>OUT_1</name></connection>
<intersection>288.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>288.5,-173,307,-173</points>
<connection>
<GID>597</GID>
<name>IN_1</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,-178.5,287.5,-145.5</points>
<intersection>-178.5 3</intersection>
<intersection>-162 2</intersection>
<intersection>-145.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287.5,-145.5,306.5,-145.5</points>
<connection>
<GID>617</GID>
<name>IN_B_0</name></connection>
<intersection>287.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-162,287.5,-162</points>
<connection>
<GID>593</GID>
<name>OUT_0</name></connection>
<intersection>287.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>287.5,-178.5,307,-178.5</points>
<connection>
<GID>598</GID>
<name>IN_1</name></connection>
<intersection>287.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-141,286,-139.5</points>
<intersection>-141 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-139.5,306.5,-139.5</points>
<connection>
<GID>616</GID>
<name>IN_3</name></connection>
<intersection>286 0</intersection>
<intersection>306 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-141,286,-141</points>
<connection>
<GID>592</GID>
<name>OUT_3</name></connection>
<intersection>286 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>306,-182,306,-139.5</points>
<intersection>-182 4</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>306,-182,307,-182</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>306 3</intersection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285,-187.5,285,-138.5</points>
<intersection>-187.5 3</intersection>
<intersection>-143 2</intersection>
<intersection>-138.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>285,-138.5,306.5,-138.5</points>
<connection>
<GID>616</GID>
<name>IN_2</name></connection>
<intersection>285 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-143,285,-143</points>
<connection>
<GID>592</GID>
<name>OUT_2</name></connection>
<intersection>285 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>285,-187.5,307,-187.5</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<intersection>285 0</intersection></hsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-192.5,284,-137.5</points>
<intersection>-192.5 3</intersection>
<intersection>-145 2</intersection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284,-137.5,306.5,-137.5</points>
<connection>
<GID>616</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-145,284,-145</points>
<connection>
<GID>592</GID>
<name>OUT_1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>284,-192.5,307,-192.5</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>284 0</intersection></hsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283,-198,283,-136.5</points>
<intersection>-198 3</intersection>
<intersection>-147 2</intersection>
<intersection>-136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>283,-136.5,306.5,-136.5</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<intersection>283 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-147,283,-147</points>
<connection>
<GID>592</GID>
<name>OUT_0</name></connection>
<intersection>283 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>283,-198,307,-198</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<intersection>283 0</intersection></hsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292.5,-184,292.5,-132.5</points>
<intersection>-184 3</intersection>
<intersection>-170.5 2</intersection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292.5,-132.5,306.5,-132.5</points>
<connection>
<GID>616</GID>
<name>IN_B_3</name></connection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-170.5,292.5,-170.5</points>
<connection>
<GID>594</GID>
<name>OUT_3</name></connection>
<intersection>292.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>292.5,-184,307,-184</points>
<connection>
<GID>599</GID>
<name>IN_1</name></connection>
<intersection>292.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-189.5,292,-131.5</points>
<intersection>-189.5 3</intersection>
<intersection>-172.5 2</intersection>
<intersection>-131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292,-131.5,306.5,-131.5</points>
<connection>
<GID>616</GID>
<name>IN_B_2</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-172.5,292,-172.5</points>
<connection>
<GID>594</GID>
<name>OUT_2</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>292,-189.5,307,-189.5</points>
<connection>
<GID>600</GID>
<name>IN_1</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,-194.5,291.5,-130.5</points>
<intersection>-194.5 3</intersection>
<intersection>-174.5 2</intersection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>291.5,-130.5,306.5,-130.5</points>
<connection>
<GID>616</GID>
<name>IN_B_1</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-174.5,291.5,-174.5</points>
<connection>
<GID>594</GID>
<name>OUT_1</name></connection>
<intersection>291.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-194.5,307,-194.5</points>
<connection>
<GID>601</GID>
<name>IN_1</name></connection>
<intersection>291.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-200,290.5,-129.5</points>
<intersection>-200 3</intersection>
<intersection>-176.5 2</intersection>
<intersection>-129.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,-129.5,306.5,-129.5</points>
<connection>
<GID>616</GID>
<name>IN_B_0</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-176.5,290.5,-176.5</points>
<connection>
<GID>594</GID>
<name>OUT_0</name></connection>
<intersection>290.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>290.5,-200,307,-200</points>
<connection>
<GID>602</GID>
<name>IN_1</name></connection>
<intersection>290.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326.5,-184.5,326.5,-133</points>
<intersection>-184.5 1</intersection>
<intersection>-133 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>326.5,-184.5,335.5,-184.5</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<intersection>326.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314.5,-133,326.5,-133</points>
<connection>
<GID>616</GID>
<name>OUT_0</name></connection>
<intersection>326.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325.5,-179.5,325.5,-134</points>
<intersection>-179.5 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>325.5,-179.5,335.5,-179.5</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<intersection>325.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314.5,-134,325.5,-134</points>
<connection>
<GID>616</GID>
<name>OUT_1</name></connection>
<intersection>325.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324.5,-174.5,324.5,-135</points>
<intersection>-174.5 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324.5,-174.5,335.5,-174.5</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<intersection>324.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314.5,-135,324.5,-135</points>
<connection>
<GID>616</GID>
<name>OUT_2</name></connection>
<intersection>324.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323.5,-169.5,323.5,-136</points>
<intersection>-169.5 1</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323.5,-169.5,335.5,-169.5</points>
<connection>
<GID>607</GID>
<name>IN_0</name></connection>
<intersection>323.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314.5,-136,323.5,-136</points>
<connection>
<GID>616</GID>
<name>OUT_3</name></connection>
<intersection>323.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322.5,-159,322.5,-149</points>
<intersection>-159 1</intersection>
<intersection>-149 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322.5,-159,335.5,-159</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>322.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314.5,-149,322.5,-149</points>
<connection>
<GID>617</GID>
<name>OUT_0</name></connection>
<intersection>322.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321.5,-154,321.5,-150</points>
<intersection>-154 1</intersection>
<intersection>-150 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321.5,-154,335.5,-154</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>321.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314.5,-150,321.5,-150</points>
<connection>
<GID>617</GID>
<name>OUT_1</name></connection>
<intersection>321.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320.5,-151,320.5,-148.5</points>
<intersection>-151 2</intersection>
<intersection>-148.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-148.5,335.5,-148.5</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>320.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314.5,-151,320.5,-151</points>
<connection>
<GID>617</GID>
<name>OUT_2</name></connection>
<intersection>320.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-152,319.5,-143</points>
<intersection>-152 2</intersection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-143,335.5,-143</points>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>319.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314.5,-152,319.5,-152</points>
<connection>
<GID>617</GID>
<name>OUT_3</name></connection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322,-182.5,322,-161</points>
<intersection>-182.5 1</intersection>
<intersection>-161 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,-182.5,335.5,-182.5</points>
<connection>
<GID>610</GID>
<name>IN_1</name></connection>
<intersection>322 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-161,322,-161</points>
<connection>
<GID>595</GID>
<name>OUT</name></connection>
<intersection>322 0</intersection></hsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321,-177.5,321,-166.5</points>
<intersection>-177.5 1</intersection>
<intersection>-166.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321,-177.5,335.5,-177.5</points>
<connection>
<GID>609</GID>
<name>IN_1</name></connection>
<intersection>321 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-166.5,321,-166.5</points>
<connection>
<GID>596</GID>
<name>OUT</name></connection>
<intersection>321 0</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320,-172.5,320,-172</points>
<intersection>-172.5 1</intersection>
<intersection>-172 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-172.5,335.5,-172.5</points>
<connection>
<GID>608</GID>
<name>IN_1</name></connection>
<intersection>320 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-172,320,-172</points>
<connection>
<GID>597</GID>
<name>OUT</name></connection>
<intersection>320 0</intersection></hsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320,-177.5,320,-167.5</points>
<intersection>-177.5 2</intersection>
<intersection>-167.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-167.5,335.5,-167.5</points>
<connection>
<GID>607</GID>
<name>IN_1</name></connection>
<intersection>320 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-177.5,320,-177.5</points>
<connection>
<GID>598</GID>
<name>OUT</name></connection>
<intersection>320 0</intersection></hsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319,-183,319,-157</points>
<intersection>-183 2</intersection>
<intersection>-157 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,-157,335.5,-157</points>
<connection>
<GID>606</GID>
<name>IN_1</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-183,319,-183</points>
<connection>
<GID>599</GID>
<name>OUT</name></connection>
<intersection>319 0</intersection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323.5,-189,323.5,-152</points>
<intersection>-189 2</intersection>
<intersection>-152 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323.5,-152,335.5,-152</points>
<connection>
<GID>605</GID>
<name>IN_1</name></connection>
<intersection>323.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-189,323.5,-189</points>
<intersection>313 3</intersection>
<intersection>323.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>313,-189,313,-188.5</points>
<connection>
<GID>600</GID>
<name>OUT</name></connection>
<intersection>-189 2</intersection></vsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324,-193.5,324,-146.5</points>
<intersection>-193.5 2</intersection>
<intersection>-146.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324,-146.5,335.5,-146.5</points>
<connection>
<GID>604</GID>
<name>IN_1</name></connection>
<intersection>324 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-193.5,324,-193.5</points>
<connection>
<GID>601</GID>
<name>OUT</name></connection>
<intersection>324 0</intersection></hsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324.5,-199,324.5,-141</points>
<intersection>-199 2</intersection>
<intersection>-141 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324.5,-141,335.5,-141</points>
<connection>
<GID>603</GID>
<name>IN_1</name></connection>
<intersection>324.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-199,324.5,-199</points>
<connection>
<GID>602</GID>
<name>OUT</name></connection>
<intersection>324.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,-181,337.5,-128.5</points>
<connection>
<GID>610</GID>
<name>SEL_0</name></connection>
<connection>
<GID>609</GID>
<name>SEL_0</name></connection>
<connection>
<GID>608</GID>
<name>SEL_0</name></connection>
<connection>
<GID>607</GID>
<name>SEL_0</name></connection>
<connection>
<GID>606</GID>
<name>SEL_0</name></connection>
<connection>
<GID>605</GID>
<name>SEL_0</name></connection>
<connection>
<GID>604</GID>
<name>SEL_0</name></connection>
<connection>
<GID>603</GID>
<name>SEL_0</name></connection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>337.5,-128.5,339,-128.5</points>
<connection>
<GID>611</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363,-159.5,363,-142</points>
<connection>
<GID>612</GID>
<name>IN_7</name></connection>
<intersection>-142 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-142,363,-142</points>
<connection>
<GID>603</GID>
<name>OUT</name></connection>
<intersection>363 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,-160.5,361.5,-147.5</points>
<intersection>-160.5 1</intersection>
<intersection>-147.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361.5,-160.5,363,-160.5</points>
<connection>
<GID>612</GID>
<name>IN_6</name></connection>
<intersection>361.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-147.5,361.5,-147.5</points>
<connection>
<GID>604</GID>
<name>OUT</name></connection>
<intersection>361.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>360,-161.5,360,-153</points>
<intersection>-161.5 1</intersection>
<intersection>-153 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,-161.5,363,-161.5</points>
<connection>
<GID>612</GID>
<name>IN_5</name></connection>
<intersection>360 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-153,360,-153</points>
<connection>
<GID>605</GID>
<name>OUT</name></connection>
<intersection>360 0</intersection></hsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-162.5,359,-158</points>
<intersection>-162.5 1</intersection>
<intersection>-158 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-162.5,363,-162.5</points>
<connection>
<GID>612</GID>
<name>IN_4</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-158,359,-158</points>
<connection>
<GID>606</GID>
<name>OUT</name></connection>
<intersection>359 0</intersection></hsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-168.5,359,-163.5</points>
<intersection>-168.5 2</intersection>
<intersection>-163.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-163.5,363,-163.5</points>
<connection>
<GID>612</GID>
<name>IN_3</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-168.5,359,-168.5</points>
<connection>
<GID>607</GID>
<name>OUT</name></connection>
<intersection>359 0</intersection></hsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>360,-173.5,360,-164.5</points>
<intersection>-173.5 2</intersection>
<intersection>-164.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,-164.5,363,-164.5</points>
<connection>
<GID>612</GID>
<name>IN_2</name></connection>
<intersection>360 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-173.5,360,-173.5</points>
<connection>
<GID>608</GID>
<name>OUT</name></connection>
<intersection>360 0</intersection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,-178.5,361.5,-165.5</points>
<intersection>-178.5 2</intersection>
<intersection>-165.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361.5,-165.5,363,-165.5</points>
<connection>
<GID>612</GID>
<name>IN_1</name></connection>
<intersection>361.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-178.5,361.5,-178.5</points>
<connection>
<GID>609</GID>
<name>OUT</name></connection>
<intersection>361.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363,-183.5,363,-166.5</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>-183.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>339.5,-183.5,363,-183.5</points>
<connection>
<GID>610</GID>
<name>OUT</name></connection>
<intersection>363 0</intersection></hsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>518.5,-128,518.5,-47.5</points>
<intersection>-128 2</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>480,-47.5,518.5,-47.5</points>
<connection>
<GID>545</GID>
<name>OUT_0</name></connection>
<intersection>518.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>518.5,-128,612,-128</points>
<connection>
<GID>571</GID>
<name>IN_2</name></connection>
<intersection>518.5 0</intersection>
<intersection>599 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>599,-128,599,-118.5</points>
<intersection>-128 2</intersection>
<intersection>-118.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>599,-118.5,605,-118.5</points>
<connection>
<GID>570</GID>
<name>IN_2</name></connection>
<intersection>599 3</intersection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>527,-126,527,-23.5</points>
<intersection>-126 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,-23.5,527,-23.5</points>
<connection>
<GID>529</GID>
<name>OUT_0</name></connection>
<intersection>527 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>527,-126,612,-126</points>
<connection>
<GID>571</GID>
<name>IN_3</name></connection>
<intersection>527 0</intersection>
<intersection>597 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>597,-126,597,-116.5</points>
<intersection>-126 2</intersection>
<intersection>-116.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>597,-116.5,605,-116.5</points>
<connection>
<GID>570</GID>
<name>IN_3</name></connection>
<intersection>597 3</intersection></hsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,-119.5,618.5,-27</points>
<intersection>-119.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,-27,650,-27</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<intersection>618.5 0</intersection>
<intersection>650 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>611,-119.5,618.5,-119.5</points>
<connection>
<GID>570</GID>
<name>OUT</name></connection>
<intersection>618.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>650,-40.5,650,-27</points>
<intersection>-40.5 4</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>650,-40.5,669,-40.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>650 3</intersection></hsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>628,-129,628,-67.5</points>
<intersection>-129 8</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>628,-67.5,652,-67.5</points>
<intersection>628 0</intersection>
<intersection>652 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>652,-79,652,-65</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>-79 5</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>652,-79,671,-79</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>652 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>618,-129,628,-129</points>
<connection>
<GID>571</GID>
<name>OUT</name></connection>
<intersection>628 0</intersection></hsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539,-112,539,-96.5</points>
<intersection>-112 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-96.5,539,-96.5</points>
<connection>
<GID>557</GID>
<name>OUT_1</name></connection>
<intersection>539 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>539,-112,598.5,-112</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>539 0</intersection>
<intersection>590 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>590,-112,590,-102</points>
<intersection>-112 2</intersection>
<intersection>-102 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>590,-102,593,-102</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>590 3</intersection></hsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539,-110,539,-71.5</points>
<intersection>-110 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>479.5,-71.5,539,-71.5</points>
<connection>
<GID>555</GID>
<name>OUT_1</name></connection>
<intersection>539 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>539,-110,598.5,-110</points>
<connection>
<GID>575</GID>
<name>IN_1</name></connection>
<intersection>539 0</intersection>
<intersection>587.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>587.5,-110,587.5,-100</points>
<intersection>-110 2</intersection>
<intersection>-100 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>587.5,-100,593,-100</points>
<connection>
<GID>574</GID>
<name>IN_1</name></connection>
<intersection>587.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539,-108,539,-46.5</points>
<intersection>-108 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>480,-46.5,539,-46.5</points>
<connection>
<GID>545</GID>
<name>OUT_1</name></connection>
<intersection>539 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>539,-108,598.5,-108</points>
<connection>
<GID>575</GID>
<name>IN_2</name></connection>
<intersection>539 0</intersection>
<intersection>585 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>585,-108,585,-98</points>
<intersection>-108 2</intersection>
<intersection>-98 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>585,-98,593,-98</points>
<connection>
<GID>574</GID>
<name>IN_2</name></connection>
<intersection>585 3</intersection></hsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539,-106,539,-22.5</points>
<intersection>-106 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,-22.5,539,-22.5</points>
<connection>
<GID>529</GID>
<name>OUT_1</name></connection>
<intersection>539 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>539,-106,598.5,-106</points>
<connection>
<GID>575</GID>
<name>IN_3</name></connection>
<intersection>539 0</intersection>
<intersection>582.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>582.5,-106,582.5,-96</points>
<intersection>-106 2</intersection>
<intersection>-96 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>582.5,-96,593,-96</points>
<connection>
<GID>574</GID>
<name>IN_3</name></connection>
<intersection>582.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>627,-109,627,-26</points>
<intersection>-109 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>627,-26,650,-26</points>
<connection>
<GID>569</GID>
<name>IN_1</name></connection>
<intersection>627 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>604.5,-109,627,-109</points>
<connection>
<GID>575</GID>
<name>OUT</name></connection>
<intersection>627 0</intersection></hsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>625.5,-99,625.5,-64</points>
<intersection>-99 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>625.5,-64,652,-64</points>
<connection>
<GID>454</GID>
<name>IN_1</name></connection>
<intersection>625.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>599,-99,625.5,-99</points>
<connection>
<GID>574</GID>
<name>OUT</name></connection>
<intersection>625.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-38,225,-19.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<connection>
<GID>644</GID>
<name>DATA_OUT_11</name></connection></vsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207.5,56,223.5,56</points>
<connection>
<GID>480</GID>
<name>OUT_4</name></connection>
<connection>
<GID>395</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,38.5,289,46</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>38.5 2</intersection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,40.5,290.5,40.5</points>
<connection>
<GID>398</GID>
<name>OUT_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>289,38.5,290.5,38.5</points>
<connection>
<GID>498</GID>
<name>count_enable</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,39.5,293.5,40.5</points>
<connection>
<GID>408</GID>
<name>OUT_0</name></connection>
<intersection>39.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>291.5,38.5,291.5,39.5</points>
<connection>
<GID>498</GID>
<name>count_up</name></connection>
<intersection>39.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>291.5,39.5,293.5,39.5</points>
<intersection>291.5 1</intersection>
<intersection>293.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,23,293,27.5</points>
<intersection>23 2</intersection>
<intersection>27.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>297.5,23,297.5,23.5</points>
<connection>
<GID>426</GID>
<name>OUT_0</name></connection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>293,23,297.5,23</points>
<intersection>293 0</intersection>
<intersection>297.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>291.5,27.5,293,27.5</points>
<connection>
<GID>498</GID>
<name>clear</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-9,237.5,11.5</points>
<connection>
<GID>644</GID>
<name>ENABLE_0</name></connection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>237.5,11.5,238,11.5</points>
<connection>
<GID>449</GID>
<name>OUT_0</name></connection>
<intersection>237.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-18.5,136,-13.5</points>
<intersection>-18.5 1</intersection>
<intersection>-13.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-18.5,136,-18.5</points>
<connection>
<GID>494</GID>
<name>ENABLE_0</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>136,-13.5,138,-13.5</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-287.367,194.69,347.872,-158.574</PageViewport></page 1>
<page 2>
<PageViewport>-11.003,20.439,689.151,-368.926</PageViewport></page 2>
<page 3>
<PageViewport>-30.9172,78.7164,839.856,-405.532</PageViewport>
<gate>
<ID>58</ID>
<type>DD_KEYPAD_HEX</type>
<position>48.5,-10.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<output>
<ID>OUT_1</ID>92 </output>
<output>
<ID>OUT_2</ID>91 </output>
<output>
<ID>OUT_3</ID>90 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_REGISTER8</type>
<position>39.5,-21.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>67 </input>
<input>
<ID>IN_2</ID>66 </input>
<input>
<ID>IN_3</ID>65 </input>
<input>
<ID>IN_4</ID>64 </input>
<input>
<ID>IN_5</ID>63 </input>
<input>
<ID>IN_6</ID>62 </input>
<input>
<ID>IN_7</ID>61 </input>
<output>
<ID>OUT_0</ID>69 </output>
<output>
<ID>OUT_1</ID>70 </output>
<output>
<ID>OUT_2</ID>71 </output>
<output>
<ID>OUT_3</ID>72 </output>
<output>
<ID>OUT_4</ID>95 </output>
<output>
<ID>OUT_5</ID>96 </output>
<output>
<ID>OUT_6</ID>97 </output>
<output>
<ID>OUT_7</ID>94 </output>
<input>
<ID>clear</ID>60 </input>
<input>
<ID>clock</ID>59 </input>
<input>
<ID>count_enable</ID>103 </input>
<input>
<ID>load</ID>102 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_REGISTER8</type>
<position>116,-55.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>67 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>66 </input>
<input>
<ID>IN_5</ID>62 </input>
<input>
<ID>IN_6</ID>65 </input>
<input>
<ID>IN_7</ID>61 </input>
<output>
<ID>OUT_0</ID>54 </output>
<output>
<ID>OUT_1</ID>53 </output>
<output>
<ID>OUT_2</ID>52 </output>
<output>
<ID>OUT_3</ID>51 </output>
<output>
<ID>OUT_4</ID>50 </output>
<output>
<ID>OUT_5</ID>49 </output>
<output>
<ID>OUT_6</ID>48 </output>
<output>
<ID>OUT_7</ID>47 </output>
<input>
<ID>clear</ID>56 </input>
<input>
<ID>clock</ID>55 </input>
<input>
<ID>load</ID>57 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_FULLADDER_4BIT</type>
<position>52.5,-33</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<input>
<ID>IN_2</ID>71 </input>
<input>
<ID>IN_3</ID>72 </input>
<input>
<ID>IN_B_0</ID>93 </input>
<input>
<ID>IN_B_1</ID>92 </input>
<input>
<ID>IN_B_2</ID>91 </input>
<input>
<ID>IN_B_3</ID>90 </input>
<output>
<ID>OUT_0</ID>89 </output>
<output>
<ID>OUT_1</ID>88 </output>
<output>
<ID>OUT_2</ID>87 </output>
<output>
<ID>OUT_3</ID>86 </output>
<output>
<ID>carry_out</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_FULLADDER_4BIT</type>
<position>69.5,-33</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>96 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>94 </input>
<input>
<ID>IN_B_0</ID>99 </input>
<input>
<ID>IN_B_1</ID>99 </input>
<input>
<ID>IN_B_2</ID>99 </input>
<input>
<ID>IN_B_3</ID>99 </input>
<output>
<ID>OUT_0</ID>81 </output>
<output>
<ID>OUT_1</ID>80 </output>
<output>
<ID>OUT_2</ID>79 </output>
<output>
<ID>OUT_3</ID>74 </output>
<input>
<ID>carry_in</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_FULLADDER_4BIT</type>
<position>88.5,-33</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<input>
<ID>IN_2</ID>71 </input>
<input>
<ID>IN_3</ID>72 </input>
<input>
<ID>IN_B_0</ID>100 </input>
<input>
<ID>IN_B_1</ID>99 </input>
<input>
<ID>IN_B_2</ID>99 </input>
<input>
<ID>IN_B_3</ID>99 </input>
<output>
<ID>OUT_0</ID>85 </output>
<output>
<ID>OUT_1</ID>84 </output>
<output>
<ID>OUT_2</ID>83 </output>
<output>
<ID>OUT_3</ID>82 </output>
<output>
<ID>carry_out</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_FULLADDER_4BIT</type>
<position>105.5,-33</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>96 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>94 </input>
<input>
<ID>IN_B_0</ID>98 </input>
<input>
<ID>IN_B_1</ID>98 </input>
<input>
<ID>IN_B_2</ID>98 </input>
<input>
<ID>IN_B_3</ID>98 </input>
<output>
<ID>OUT_0</ID>78 </output>
<output>
<ID>OUT_1</ID>77 </output>
<output>
<ID>OUT_2</ID>76 </output>
<output>
<ID>OUT_3</ID>75 </output>
<input>
<ID>carry_in</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>65</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>123,-55</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>53 </input>
<input>
<ID>IN_2</ID>52 </input>
<input>
<ID>IN_3</ID>51 </input>
<input>
<ID>IN_4</ID>50 </input>
<input>
<ID>IN_5</ID>49 </input>
<input>
<ID>IN_6</ID>48 </input>
<input>
<ID>IN_7</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>115,-46.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>117,-63.5</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>40.5,-29.5</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_TOGGLE</type>
<position>35.5,-14</position>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_TOGGLE</type>
<position>35.5,-11</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>49.5,-80</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>72</ID>
<type>FF_GND</type>
<position>109,-26</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>FF_GND</type>
<position>73,-26</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>EE_VDD</type>
<position>93.5,-27</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>75</ID>
<type>BB_CLOCK</type>
<position>38.5,-34.5</position>
<output>
<ID>CLK</ID>59 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>76</ID>
<type>BB_CLOCK</type>
<position>115,-68.5</position>
<output>
<ID>CLK</ID>55 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_MUX_2x1</type>
<position>45,-54.5</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>66 </output>
<input>
<ID>SEL_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_MUX_2x1</type>
<position>60,-49</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>62 </output>
<input>
<ID>SEL_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_MUX_2x1</type>
<position>42,-45.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>65 </output>
<input>
<ID>SEL_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_MUX_2x1</type>
<position>48,-64.5</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>67 </output>
<input>
<ID>SEL_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_MUX_2x1</type>
<position>57,-41</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>61 </output>
<input>
<ID>SEL_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_MUX_2x1</type>
<position>63,-59</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>63 </output>
<input>
<ID>SEL_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_MUX_2x1</type>
<position>51,-73.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>68 </output>
<input>
<ID>SEL_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_MUX_2x1</type>
<position>66,-68</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>64 </output>
<input>
<ID>SEL_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>48.5,-2</position>
<gparam>LABEL_TEXT PCOffset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>27,-10.5</position>
<gparam>LABEL_TEXT Countup</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>29.5,-13.5</position>
<gparam>LABEL_TEXT Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>44,-27.5</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>134.5,-54.5</position>
<gparam>LABEL_TEXT Global Bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>123.5,-63</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>115,-43</position>
<gparam>LABEL_TEXT Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>49.5,-82.5</position>
<gparam>LABEL_TEXT Most/Least Significant</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>120,-51.5,121,-51.5</points>
<connection>
<GID>60</GID>
<name>OUT_7</name></connection>
<connection>
<GID>65</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>120,-52.5,121,-52.5</points>
<connection>
<GID>60</GID>
<name>OUT_6</name></connection>
<connection>
<GID>65</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>120,-53.5,121,-53.5</points>
<connection>
<GID>60</GID>
<name>OUT_5</name></connection>
<connection>
<GID>65</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>120,-54.5,121,-54.5</points>
<connection>
<GID>60</GID>
<name>OUT_4</name></connection>
<connection>
<GID>65</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>120,-55.5,121,-55.5</points>
<connection>
<GID>60</GID>
<name>OUT_3</name></connection>
<connection>
<GID>65</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>120,-56.5,121,-56.5</points>
<connection>
<GID>60</GID>
<name>OUT_2</name></connection>
<connection>
<GID>65</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>120,-57.5,121,-57.5</points>
<connection>
<GID>60</GID>
<name>OUT_1</name></connection>
<connection>
<GID>65</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>120,-58.5,121,-58.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>20</ID>
<points>115,-64.5,115,-60.5</points>
<connection>
<GID>76</GID>
<name>CLK</name></connection>
<connection>
<GID>60</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>117,-61.5,117,-60.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<connection>
<GID>60</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>26</ID>
<points>115,-49.5,115,-48.5</points>
<connection>
<GID>60</GID>
<name>load</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,-38,78.5,-38</points>
<intersection>43.5 7</intersection>
<intersection>78.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>78.5,-38,78.5,-32</points>
<intersection>-38 1</intersection>
<intersection>-32 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>77.5,-32,78.5,-32</points>
<connection>
<GID>62</GID>
<name>carry_in</name></connection>
<intersection>78.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>43.5,-38,43.5,-32</points>
<intersection>-38 1</intersection>
<intersection>-32 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>43.5,-32,44.5,-32</points>
<connection>
<GID>61</GID>
<name>carry_out</name></connection>
<intersection>43.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>38.5,-30.5,38.5,-26.5</points>
<connection>
<GID>75</GID>
<name>CLK</name></connection>
<connection>
<GID>59</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>40.5,-27.5,40.5,-26.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-41,110,-41</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<intersection>34.5 3</intersection>
<intersection>110 10</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34.5,-41,34.5,-17.5</points>
<intersection>-41 1</intersection>
<intersection>-17.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>34.5,-17.5,35.5,-17.5</points>
<connection>
<GID>59</GID>
<name>IN_7</name></connection>
<intersection>34.5 3</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>110,-51.5,110,-41</points>
<intersection>-51.5 11</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>110,-51.5,112,-51.5</points>
<connection>
<GID>60</GID>
<name>IN_7</name></connection>
<intersection>110 10</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-49,33.5,-18.5</points>
<intersection>-49 1</intersection>
<intersection>-18.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-49,108,-49</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>33.5 0</intersection>
<intersection>108 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-18.5,35.5,-18.5</points>
<connection>
<GID>59</GID>
<name>IN_6</name></connection>
<intersection>33.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>108,-53.5,108,-49</points>
<intersection>-53.5 5</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>108,-53.5,112,-53.5</points>
<connection>
<GID>60</GID>
<name>IN_5</name></connection>
<intersection>108 4</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-59,32.5,-19.5</points>
<intersection>-59 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-59,108,-59</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection>
<intersection>108 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-19.5,35.5,-19.5</points>
<connection>
<GID>59</GID>
<name>IN_5</name></connection>
<intersection>32.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>108,-59,108,-55.5</points>
<intersection>-59 1</intersection>
<intersection>-55.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>108,-55.5,112,-55.5</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>108 3</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-68,31.5,-20.5</points>
<intersection>-68 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-20.5,35.5,-20.5</points>
<connection>
<GID>59</GID>
<name>IN_4</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-68,110,-68</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<intersection>31.5 0</intersection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,-68,110,-57.5</points>
<intersection>-68 2</intersection>
<intersection>-57.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>110,-57.5,112,-57.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>110 3</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-45.5,30.5,-21.5</points>
<intersection>-45.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-45.5,109,-45.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>30.5 0</intersection>
<intersection>109 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-21.5,35.5,-21.5</points>
<connection>
<GID>59</GID>
<name>IN_3</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109,-52.5,109,-45.5</points>
<intersection>-52.5 4</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>109,-52.5,112,-52.5</points>
<connection>
<GID>60</GID>
<name>IN_6</name></connection>
<intersection>109 3</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-54.5,29.5,-22.5</points>
<intersection>-54.5 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-54.5,112,-54.5</points>
<connection>
<GID>60</GID>
<name>IN_4</name></connection>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-22.5,35.5,-22.5</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-64.5,28.5,-23.5</points>
<intersection>-64.5 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-64.5,109,-64.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection>
<intersection>109 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-23.5,35.5,-23.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109,-64.5,109,-56.5</points>
<intersection>-64.5 1</intersection>
<intersection>-56.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>109,-56.5,112,-56.5</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>109 3</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-73.5,27.5,-24.5</points>
<intersection>-73.5 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-73.5,111,-73.5</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection>
<intersection>111 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-24.5,35.5,-24.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111,-73.5,111,-58.5</points>
<intersection>-73.5 1</intersection>
<intersection>-58.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>111,-58.5,112,-58.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>111 3</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,-24.5,86.5,-24.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>50.5 5</intersection>
<intersection>86.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>86.5,-29,86.5,-24.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>50.5,-29,50.5,-24.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-29,49.5,-23.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-23.5,85.5,-23.5</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<intersection>49.5 0</intersection>
<intersection>85.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>85.5,-29,85.5,-23.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-29,48.5,-22.5</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-22.5,84.5,-22.5</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<intersection>48.5 0</intersection>
<intersection>84.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>84.5,-29,84.5,-22.5</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<intersection>-22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-29,47.5,-21.5</points>
<connection>
<GID>61</GID>
<name>IN_3</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-21.5,83.5,-21.5</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<intersection>47.5 0</intersection>
<intersection>83.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83.5,-29,83.5,-21.5</points>
<connection>
<GID>63</GID>
<name>IN_3</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,-38,114.5,-38</points>
<intersection>79.5 4</intersection>
<intersection>114.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114.5,-38,114.5,-32</points>
<intersection>-38 1</intersection>
<intersection>-32 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>79.5,-38,79.5,-32</points>
<intersection>-38 1</intersection>
<intersection>-32 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>79.5,-32,80.5,-32</points>
<connection>
<GID>63</GID>
<name>carry_out</name></connection>
<intersection>79.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>113.5,-32,114.5,-32</points>
<connection>
<GID>64</GID>
<name>carry_in</name></connection>
<intersection>114.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-42,68,-37</points>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-42,68,-42</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-40,104,-37</points>
<connection>
<GID>64</GID>
<name>OUT_3</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-40,104,-40</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-48,105,-37</points>
<connection>
<GID>64</GID>
<name>OUT_2</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-48,105,-48</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-58,106,-37</points>
<connection>
<GID>64</GID>
<name>OUT_1</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-58,106,-58</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-67,107,-37</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-67,107,-67</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-50,69,-37</points>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-50,69,-50</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-60,70,-37</points>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-60,70,-60</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-69,71,-37</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-69,71,-69</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-44.5,87,-37</points>
<connection>
<GID>63</GID>
<name>OUT_3</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-44.5,87,-44.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-53.5,88,-37</points>
<connection>
<GID>63</GID>
<name>OUT_2</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-53.5,88,-53.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-63.5,89,-37</points>
<connection>
<GID>63</GID>
<name>OUT_1</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-63.5,89,-63.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-72.5,90,-37</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-72.5,90,-72.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-46.5,51,-37</points>
<connection>
<GID>61</GID>
<name>OUT_3</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-46.5,51,-46.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-55.5,52,-37</points>
<connection>
<GID>61</GID>
<name>OUT_2</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-55.5,52,-55.5</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-65.5,53,-37</points>
<connection>
<GID>61</GID>
<name>OUT_1</name></connection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-65.5,53,-65.5</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-74.5,54,-37</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-74.5,54,-74.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-29,54.5,-7.5</points>
<connection>
<GID>61</GID>
<name>IN_B_3</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-7.5,54.5,-7.5</points>
<connection>
<GID>58</GID>
<name>OUT_3</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-29,55.5,-9.5</points>
<connection>
<GID>61</GID>
<name>IN_B_2</name></connection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-9.5,55.5,-9.5</points>
<connection>
<GID>58</GID>
<name>OUT_2</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-29,56.5,-11.5</points>
<connection>
<GID>61</GID>
<name>IN_B_1</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-11.5,56.5,-11.5</points>
<connection>
<GID>58</GID>
<name>OUT_1</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-29,57.5,-13.5</points>
<connection>
<GID>61</GID>
<name>IN_B_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-13.5,57.5,-13.5</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-29,64.5,-17.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-17.5,100.5,-17.5</points>
<connection>
<GID>59</GID>
<name>OUT_7</name></connection>
<intersection>64.5 0</intersection>
<intersection>100.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100.5,-29,100.5,-17.5</points>
<connection>
<GID>64</GID>
<name>IN_3</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-29,67.5,-20.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-20.5,103.5,-20.5</points>
<connection>
<GID>59</GID>
<name>OUT_4</name></connection>
<intersection>67.5 0</intersection>
<intersection>103.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>103.5,-29,103.5,-20.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-29,66.5,-19.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-19.5,102.5,-19.5</points>
<connection>
<GID>59</GID>
<name>OUT_5</name></connection>
<intersection>66.5 0</intersection>
<intersection>102.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>102.5,-29,102.5,-19.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>-19.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-29,65.5,-18.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-18.5,101.5,-18.5</points>
<connection>
<GID>59</GID>
<name>OUT_6</name></connection>
<intersection>65.5 0</intersection>
<intersection>101.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>101.5,-29,101.5,-18.5</points>
<connection>
<GID>64</GID>
<name>IN_2</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-29,109.5,-28</points>
<connection>
<GID>64</GID>
<name>IN_B_1</name></connection>
<intersection>-28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107.5,-28,110.5,-28</points>
<intersection>107.5 4</intersection>
<intersection>108.5 5</intersection>
<intersection>109 12</intersection>
<intersection>109.5 0</intersection>
<intersection>110.5 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>107.5,-29,107.5,-28</points>
<connection>
<GID>64</GID>
<name>IN_B_3</name></connection>
<intersection>-28 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>108.5,-29,108.5,-28</points>
<connection>
<GID>64</GID>
<name>IN_B_2</name></connection>
<intersection>-28 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>110.5,-29,110.5,-28</points>
<connection>
<GID>64</GID>
<name>IN_B_0</name></connection>
<intersection>-28 3</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>109,-28,109,-27</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-28 3</intersection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-29,71.5,-28</points>
<connection>
<GID>62</GID>
<name>IN_B_3</name></connection>
<intersection>-28 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>71.5,-28,92.5,-28</points>
<intersection>71.5 0</intersection>
<intersection>72.5 6</intersection>
<intersection>73 4</intersection>
<intersection>73.5 8</intersection>
<intersection>74.5 10</intersection>
<intersection>90.5 12</intersection>
<intersection>91.5 14</intersection>
<intersection>92.5 16</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>73,-28,73,-27</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>-28 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>72.5,-29,72.5,-28</points>
<connection>
<GID>62</GID>
<name>IN_B_2</name></connection>
<intersection>-28 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>73.5,-29,73.5,-28</points>
<connection>
<GID>62</GID>
<name>IN_B_1</name></connection>
<intersection>-28 3</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>74.5,-29,74.5,-28</points>
<connection>
<GID>62</GID>
<name>IN_B_0</name></connection>
<intersection>-28 3</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>90.5,-29,90.5,-28</points>
<connection>
<GID>63</GID>
<name>IN_B_3</name></connection>
<intersection>-28 3</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>91.5,-29,91.5,-28</points>
<connection>
<GID>63</GID>
<name>IN_B_2</name></connection>
<intersection>-28 3</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>92.5,-29,92.5,-28</points>
<connection>
<GID>63</GID>
<name>IN_B_1</name></connection>
<intersection>-28 3</intersection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>93.5,-29,93.5,-28</points>
<connection>
<GID>63</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>42,-77,42,-48</points>
<connection>
<GID>79</GID>
<name>SEL_0</name></connection>
<intersection>-77 2</intersection>
<intersection>-67 4</intersection>
<intersection>-58 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42,-77,57,-77</points>
<intersection>42 1</intersection>
<intersection>49.5 23</intersection>
<intersection>51 27</intersection>
<intersection>57 7</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>42,-58,45,-58</points>
<intersection>42 1</intersection>
<intersection>45 15</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>42,-67,48,-67</points>
<connection>
<GID>80</GID>
<name>SEL_0</name></connection>
<intersection>42 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>57,-77,57,-43.5</points>
<connection>
<GID>81</GID>
<name>SEL_0</name></connection>
<intersection>-77 2</intersection>
<intersection>-71.5 14</intersection>
<intersection>-62.5 11</intersection>
<intersection>-52.5 13</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>57,-62.5,63,-62.5</points>
<intersection>57 7</intersection>
<intersection>63 20</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>57,-52.5,60,-52.5</points>
<intersection>57 7</intersection>
<intersection>60 16</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>57,-71.5,66,-71.5</points>
<intersection>57 7</intersection>
<intersection>66 22</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>45,-58,45,-57</points>
<connection>
<GID>77</GID>
<name>SEL_0</name></connection>
<intersection>-58 3</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>60,-52.5,60,-51.5</points>
<connection>
<GID>78</GID>
<name>SEL_0</name></connection>
<intersection>-52.5 13</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>63,-62.5,63,-61.5</points>
<connection>
<GID>82</GID>
<name>SEL_0</name></connection>
<intersection>-62.5 11</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>66,-71.5,66,-70.5</points>
<connection>
<GID>84</GID>
<name>SEL_0</name></connection>
<intersection>-71.5 14</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>49.5,-78,49.5,-77</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>-77 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>51,-77,51,-76</points>
<connection>
<GID>83</GID>
<name>SEL_0</name></connection>
<intersection>-77 2</intersection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-15.5,38.5,-14</points>
<connection>
<GID>59</GID>
<name>load</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-14,38.5,-14</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-15.5,39.5,-11</points>
<connection>
<GID>59</GID>
<name>count_enable</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-11,39.5,-11</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-324.985,234.045,640.615,-302.937</PageViewport>
<gate>
<ID>390</ID>
<type>DE_TO</type>
<position>36,29</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRload</lparam></gate>
<gate>
<ID>392</ID>
<type>DE_TO</type>
<position>36.5,33.5</position>
<input>
<ID>IN_0</ID>357 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRsend</lparam></gate>
<gate>
<ID>393</ID>
<type>DA_FROM</type>
<position>-1,146</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRrecieve</lparam></gate>
<gate>
<ID>4</ID>
<type>DD_KEYPAD_HEX</type>
<position>-112.5,-30.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>-103.5,-26</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 0</lparam></gate>
<gate>
<ID>6</ID>
<type>DE_TO</type>
<position>-103.5,-29</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 1</lparam></gate>
<gate>
<ID>7</ID>
<type>DE_TO</type>
<position>-103.5,-32</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 2</lparam></gate>
<gate>
<ID>8</ID>
<type>DE_TO</type>
<position>-103.5,-35</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 3</lparam></gate>
<gate>
<ID>9</ID>
<type>DE_TO</type>
<position>-103.5,-38</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 4</lparam></gate>
<gate>
<ID>10</ID>
<type>DE_TO</type>
<position>-103.5,-41</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 5</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>-103.5,-44</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 6</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>-103.5,-47</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SExt 7</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>21.5,-73.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-3.5,-42.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>19 </input>
<input>
<ID>IN_3</ID>20 </input>
<input>
<ID>IN_B_0</ID>16 </input>
<input>
<ID>IN_B_1</ID>15 </input>
<input>
<ID>IN_B_2</ID>14 </input>
<input>
<ID>IN_B_3</ID>13 </input>
<output>
<ID>OUT_0</ID>23 </output>
<output>
<ID>OUT_1</ID>22 </output>
<output>
<ID>OUT_2</ID>21 </output>
<output>
<ID>OUT_3</ID>29 </output>
<output>
<ID>carry_out</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>15</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-57.5,-42.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>8 </input>
<input>
<ID>IN_B_0</ID>9 </input>
<input>
<ID>IN_B_1</ID>10 </input>
<input>
<ID>IN_B_2</ID>11 </input>
<input>
<ID>IN_B_3</ID>12 </input>
<output>
<ID>OUT_0</ID>35 </output>
<output>
<ID>OUT_1</ID>37 </output>
<output>
<ID>OUT_2</ID>38 </output>
<output>
<ID>OUT_3</ID>39 </output>
<input>
<ID>carry_in</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>405</ID>
<type>DE_TO</type>
<position>37.5,37.5</position>
<input>
<ID>IN_0</ID>442 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRrecieve</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_MUX_2x1</type>
<position>-11,-58.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>31 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_MUX_2x1</type>
<position>-38,-64.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>407</ID>
<type>DA_FROM</type>
<position>196,-23.5</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load bit 4 (DR)</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_MUX_2x1</type>
<position>-51.5,-67.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>43 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_MUX_2x1</type>
<position>16,-52.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>26 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>DE_TO</type>
<position>36,131.5</position>
<input>
<ID>IN_0</ID>443 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load bit 4 (DR)</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_MUX_2x1</type>
<position>-78.5,-73.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>45 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_MUX_2x1</type>
<position>-24.5,-61.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>32 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>AA_TOGGLE</type>
<position>101,118</position>
<output>
<ID>OUT_0</ID>444 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_MUX_2x1</type>
<position>-65,-70.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>44 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_MUX_2x1</type>
<position>2,-55.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>28 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>-50,-32.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt5</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>1,-32.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt2</lparam></gate>
<gate>
<ID>415</ID>
<type>AA_TOGGLE</type>
<position>104,118</position>
<output>
<ID>OUT_0</ID>445 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>-47,-32.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt4</lparam></gate>
<gate>
<ID>27</ID>
<type>DA_FROM</type>
<position>-82.5,-48.5</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp7</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>-55.5,-50.5</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp5</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>-42,-49.5</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp4</lparam></gate>
<gate>
<ID>419</ID>
<type>DA_FROM</type>
<position>96.5,126.5</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Load</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>-5,-32.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut0</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>4,-32.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt1</lparam></gate>
<gate>
<ID>421</ID>
<type>DA_FROM</type>
<position>99.5,123.5</position>
<input>
<ID>IN_0</ID>444 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID CEnable</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>12,-49.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID PCUp0</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>-2,-32.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt3</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>-53,-32.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt6</lparam></gate>
<gate>
<ID>424</ID>
<type>AA_TOGGLE</type>
<position>108,101</position>
<output>
<ID>OUT_0</ID>446 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>7,-32.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt0</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>-1.5,-50.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID PCUp1</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>-15,-49.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID PCUp2</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>-69,-49.5</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp6</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>-28.5,-48.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCUp3</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>-11,-78.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux2</lparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>-24.5,-78.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux3</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>-38,-78.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux4</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>-78.5,-78.5</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux7</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>16,-78.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux0</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>2,-78.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux1</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>-65,-78.5</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux6</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>-51.5,-78.5</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCMux5</lparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>-56,-32.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID SExt7</lparam></gate>
<gate>
<ID>49</ID>
<type>DA_FROM</type>
<position>-11,-32.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut2</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>-59,-32.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut4</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>-65,-32.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut6</lparam></gate>
<gate>
<ID>52</ID>
<type>DA_FROM</type>
<position>-14,-32.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut3</lparam></gate>
<gate>
<ID>53</ID>
<type>DA_FROM</type>
<position>-62,-32.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut5</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>-68,-32.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut7</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>-8,-32.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCOut1</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>176,20</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>50.5,87</position>
<output>
<ID>OUT_0</ID>447 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>95</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>187.5,39</position>
<input>
<ID>ENABLE_0</ID>376 </input>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>107 </input>
<input>
<ID>IN_2</ID>108 </input>
<input>
<ID>IN_3</ID>109 </input>
<input>
<ID>IN_4</ID>112 </input>
<input>
<ID>IN_5</ID>113 </input>
<input>
<ID>IN_6</ID>114 </input>
<input>
<ID>IN_7</ID>115 </input>
<output>
<ID>OUT_0</ID>324 </output>
<output>
<ID>OUT_1</ID>323 </output>
<output>
<ID>OUT_2</ID>322 </output>
<output>
<ID>OUT_3</ID>321 </output>
<output>
<ID>OUT_4</ID>320 </output>
<output>
<ID>OUT_5</ID>319 </output>
<output>
<ID>OUT_6</ID>289 </output>
<output>
<ID>OUT_7</ID>333 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>176.5,28</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>97</ID>
<type>DA_FROM</type>
<position>174,33</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>330,137</position>
<gparam>LABEL_TEXT Register File</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>467.5,13.5</position>
<input>
<ID>IN_0</ID>435 </input>
<input>
<ID>IN_1</ID>441 </input>
<input>
<ID>IN_2</ID>134 </input>
<input>
<ID>IN_3</ID>132 </input>
<input>
<ID>IN_4</ID>130 </input>
<input>
<ID>IN_5</ID>128 </input>
<input>
<ID>IN_6</ID>361 </input>
<input>
<ID>IN_7</ID>334 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>481,58</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x7</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>480.5,51</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x5</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>480.5,48</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>480.5,44.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>481,41.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>481,38.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>481.5,35</position>
<input>
<ID>IN_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x0</lparam></gate>
<gate>
<ID>109</ID>
<type>DE_TO</type>
<position>480.5,54</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x6</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>483,20</position>
<input>
<ID>IN_0</ID>334 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y7</lparam></gate>
<gate>
<ID>111</ID>
<type>DA_FROM</type>
<position>172,38.5</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>112</ID>
<type>DA_FROM</type>
<position>155,42.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>113</ID>
<type>DA_FROM</type>
<position>156,48</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>114</ID>
<type>DA_FROM</type>
<position>155.5,52</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>115</ID>
<type>DA_FROM</type>
<position>155.5,56</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>116</ID>
<type>DE_TO</type>
<position>483.5,-3.5</position>
<input>
<ID>IN_0</ID>435 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y0</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_REGISTER8</type>
<position>-45.5,44.5</position>
<input>
<ID>IN_0</ID>232 </input>
<input>
<ID>IN_1</ID>233 </input>
<input>
<ID>IN_2</ID>234 </input>
<input>
<ID>IN_3</ID>235 </input>
<input>
<ID>IN_4</ID>278 </input>
<input>
<ID>IN_5</ID>279 </input>
<input>
<ID>IN_6</ID>280 </input>
<input>
<ID>IN_7</ID>281 </input>
<output>
<ID>OUT_0</ID>162 </output>
<output>
<ID>OUT_1</ID>161 </output>
<output>
<ID>OUT_2</ID>125 </output>
<output>
<ID>OUT_3</ID>124 </output>
<output>
<ID>OUT_4</ID>123 </output>
<output>
<ID>OUT_5</ID>122 </output>
<output>
<ID>OUT_6</ID>121 </output>
<output>
<ID>OUT_7</ID>120 </output>
<input>
<ID>clear</ID>118 </input>
<input>
<ID>clock</ID>335 </input>
<input>
<ID>load</ID>163 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>120</ID>
<type>DE_TO</type>
<position>483,17</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y6</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>112.5,161</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>-38,-14.5</position>
<gparam>LABEL_TEXT PC adder for offset in Branch Case</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>DE_TO</type>
<position>483,13</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y5</lparam></gate>
<gate>
<ID>124</ID>
<type>DE_TO</type>
<position>483,9</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y4</lparam></gate>
<gate>
<ID>125</ID>
<type>DE_TO</type>
<position>484,0</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y1</lparam></gate>
<gate>
<ID>126</ID>
<type>DE_TO</type>
<position>483.5,5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y3</lparam></gate>
<gate>
<ID>127</ID>
<type>DE_TO</type>
<position>484,2.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID y2</lparam></gate>
<gate>
<ID>128</ID>
<type>AE_REGISTER8</type>
<position>9,130.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>331 </input>
<input>
<ID>IN_2</ID>330 </input>
<input>
<ID>IN_3</ID>329 </input>
<input>
<ID>IN_4</ID>328 </input>
<input>
<ID>IN_5</ID>327 </input>
<input>
<ID>IN_6</ID>326 </input>
<input>
<ID>IN_7</ID>325 </input>
<output>
<ID>OUT_0</ID>182 </output>
<output>
<ID>OUT_1</ID>181 </output>
<output>
<ID>OUT_2</ID>180 </output>
<output>
<ID>OUT_3</ID>179 </output>
<output>
<ID>OUT_4</ID>178 </output>
<output>
<ID>OUT_5</ID>177 </output>
<output>
<ID>OUT_6</ID>176 </output>
<output>
<ID>OUT_7</ID>175 </output>
<input>
<ID>clear</ID>184 </input>
<input>
<ID>clock</ID>335 </input>
<input>
<ID>load</ID>185 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>129</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>16,131</position>
<input>
<ID>ENABLE_0</ID>366 </input>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>181 </input>
<input>
<ID>IN_2</ID>180 </input>
<input>
<ID>IN_3</ID>179 </input>
<input>
<ID>IN_4</ID>178 </input>
<input>
<ID>IN_5</ID>177 </input>
<input>
<ID>IN_6</ID>176 </input>
<input>
<ID>IN_7</ID>175 </input>
<output>
<ID>OUT_0</ID>368 </output>
<output>
<ID>OUT_1</ID>369 </output>
<output>
<ID>OUT_2</ID>370 </output>
<output>
<ID>OUT_3</ID>371 </output>
<output>
<ID>OUT_4</ID>443 </output>
<output>
<ID>OUT_5</ID>353 </output>
<output>
<ID>OUT_6</ID>364 </output>
<output>
<ID>OUT_7</ID>365 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_TOGGLE</type>
<position>10,119.5</position>
<output>
<ID>OUT_0</ID>184 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_TOGGLE</type>
<position>225.5,106</position>
<output>
<ID>OUT_0</ID>287 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>15.5,120</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>7.5,146.5</position>
<gparam>LABEL_TEXT Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>225.5,110.5</position>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>21.5,146.5</position>
<gparam>LABEL_TEXT IR control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>17.5,152</position>
<gparam>LABEL_TEXT Instruction Register</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_TOGGLE</type>
<position>-46.5,36</position>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>-46,33.5</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>466.5,61.5</position>
<gparam>LABEL_TEXT SR1 Out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_TOGGLE</type>
<position>224,121</position>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>467.5,24.5</position>
<gparam>LABEL_TEXT SR2 Out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>AA_LABEL</type>
<position>-71.5,77.5</position>
<gparam>LABEL_TEXT Memory</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>AE_RAM_8x8</type>
<position>-63,57.5</position>
<input>
<ID>ADDRESS_0</ID>202 </input>
<input>
<ID>ADDRESS_1</ID>201 </input>
<input>
<ID>ADDRESS_2</ID>200 </input>
<input>
<ID>ADDRESS_3</ID>199 </input>
<input>
<ID>ADDRESS_4</ID>198 </input>
<input>
<ID>ADDRESS_5</ID>197 </input>
<input>
<ID>ADDRESS_6</ID>196 </input>
<input>
<ID>ADDRESS_7</ID>195 </input>
<input>
<ID>DATA_IN_0</ID>232 </input>
<input>
<ID>DATA_IN_1</ID>233 </input>
<input>
<ID>DATA_IN_2</ID>234 </input>
<input>
<ID>DATA_IN_3</ID>235 </input>
<input>
<ID>DATA_IN_4</ID>278 </input>
<input>
<ID>DATA_IN_5</ID>279 </input>
<input>
<ID>DATA_IN_6</ID>280 </input>
<input>
<ID>DATA_IN_7</ID>281 </input>
<output>
<ID>DATA_OUT_0</ID>232 </output>
<output>
<ID>DATA_OUT_1</ID>233 </output>
<output>
<ID>DATA_OUT_2</ID>234 </output>
<output>
<ID>DATA_OUT_3</ID>235 </output>
<output>
<ID>DATA_OUT_4</ID>278 </output>
<output>
<ID>DATA_OUT_5</ID>279 </output>
<output>
<ID>DATA_OUT_6</ID>280 </output>
<output>
<ID>DATA_OUT_7</ID>281 </output>
<input>
<ID>ENABLE_0</ID>449 </input>
<input>
<ID>write_clock</ID>335 </input>
<input>
<ID>write_enable</ID>283 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:1 10</lparam>
<lparam>Address:2 32</lparam>
<lparam>Address:3 48</lparam>
<lparam>Address:4 64</lparam>
<lparam>Address:5 80</lparam>
<lparam>Address:6 96</lparam>
<lparam>Address:7 112</lparam></gate>
<gate>
<ID>148</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-32,45</position>
<input>
<ID>ENABLE_0</ID>119 </input>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>161 </input>
<input>
<ID>IN_2</ID>125 </input>
<input>
<ID>IN_3</ID>124 </input>
<input>
<ID>IN_4</ID>123 </input>
<input>
<ID>IN_5</ID>122 </input>
<input>
<ID>IN_6</ID>121 </input>
<input>
<ID>IN_7</ID>120 </input>
<output>
<ID>OUT_0</ID>300 </output>
<output>
<ID>OUT_1</ID>299 </output>
<output>
<ID>OUT_2</ID>298 </output>
<output>
<ID>OUT_3</ID>297 </output>
<output>
<ID>OUT_4</ID>296 </output>
<output>
<ID>OUT_5</ID>295 </output>
<output>
<ID>OUT_6</ID>294 </output>
<output>
<ID>OUT_7</ID>293 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>151</ID>
<type>DA_FROM</type>
<position>-46,53</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRload</lparam></gate>
<gate>
<ID>152</ID>
<type>DA_FROM</type>
<position>-29,52.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID MDRsend</lparam></gate>
<gate>
<ID>154</ID>
<type>AE_REGISTER8</type>
<position>101,108</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_2</ID>208 </input>
<input>
<ID>IN_3</ID>207 </input>
<input>
<ID>IN_4</ID>206 </input>
<input>
<ID>IN_5</ID>205 </input>
<input>
<ID>IN_6</ID>204 </input>
<input>
<ID>IN_7</ID>203 </input>
<output>
<ID>OUT_0</ID>218 </output>
<output>
<ID>OUT_1</ID>219 </output>
<output>
<ID>OUT_2</ID>220 </output>
<output>
<ID>OUT_3</ID>217 </output>
<output>
<ID>OUT_4</ID>213 </output>
<output>
<ID>OUT_5</ID>214 </output>
<output>
<ID>OUT_6</ID>215 </output>
<output>
<ID>OUT_7</ID>216 </output>
<input>
<ID>clear</ID>446 </input>
<input>
<ID>clock</ID>335 </input>
<input>
<ID>count_enable</ID>444 </input>
<input>
<ID>count_up</ID>445 </input>
<input>
<ID>load</ID>211 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>88.5,137</position>
<gparam>LABEL_TEXT CountIn</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>93,136.5</position>
<output>
<ID>OUT_0</ID>222 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_TOGGLE</type>
<position>98,118</position>
<output>
<ID>OUT_0</ID>211 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>90,119</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux7</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>90,116</position>
<input>
<ID>IN_0</ID>204 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux6</lparam></gate>
<gate>
<ID>161</ID>
<type>DA_FROM</type>
<position>90,113</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux5</lparam></gate>
<gate>
<ID>162</ID>
<type>DA_FROM</type>
<position>90,110</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux4</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>90,107</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux3</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>90,104</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux2</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>90,101</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux1</lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>90,98</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCMux0</lparam></gate>
<gate>
<ID>167</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>129,108.5</position>
<input>
<ID>ENABLE_0</ID>344 </input>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_2</ID>220 </input>
<input>
<ID>IN_3</ID>217 </input>
<input>
<ID>IN_4</ID>213 </input>
<input>
<ID>IN_5</ID>214 </input>
<input>
<ID>IN_6</ID>215 </input>
<input>
<ID>IN_7</ID>216 </input>
<output>
<ID>OUT_0</ID>342 </output>
<output>
<ID>OUT_1</ID>343 </output>
<output>
<ID>OUT_2</ID>345 </output>
<output>
<ID>OUT_3</ID>346 </output>
<output>
<ID>OUT_4</ID>347 </output>
<output>
<ID>OUT_5</ID>348 </output>
<output>
<ID>OUT_6</ID>349 </output>
<output>
<ID>OUT_7</ID>350 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>119.5,146.5</position>
<input>
<ID>IN_0</ID>228 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp1</lparam></gate>
<gate>
<ID>169</ID>
<type>DE_TO</type>
<position>122.5,146.5</position>
<input>
<ID>IN_0</ID>229 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp2</lparam></gate>
<gate>
<ID>170</ID>
<type>DE_TO</type>
<position>125.5,146.5</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp3</lparam></gate>
<gate>
<ID>171</ID>
<type>DE_TO</type>
<position>99.5,146.5</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp4</lparam></gate>
<gate>
<ID>172</ID>
<type>DE_TO</type>
<position>116.5,146.5</position>
<input>
<ID>IN_0</ID>231 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp0</lparam></gate>
<gate>
<ID>173</ID>
<type>DE_TO</type>
<position>102.5,146.5</position>
<input>
<ID>IN_0</ID>225 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp5</lparam></gate>
<gate>
<ID>174</ID>
<type>DE_TO</type>
<position>108.5,146.5</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp7</lparam></gate>
<gate>
<ID>175</ID>
<type>DE_TO</type>
<position>105.5,146.5</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID PCUp6</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_TOGGLE</type>
<position>224.5,124.5</position>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>177</ID>
<type>AE_FULLADDER_4BIT</type>
<position>104,137.5</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>214 </input>
<input>
<ID>IN_2</ID>215 </input>
<input>
<ID>IN_3</ID>216 </input>
<output>
<ID>OUT_0</ID>224 </output>
<output>
<ID>OUT_1</ID>225 </output>
<output>
<ID>OUT_2</ID>226 </output>
<output>
<ID>OUT_3</ID>227 </output>
<input>
<ID>carry_in</ID>222 </input>
<output>
<ID>carry_out</ID>221 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>178</ID>
<type>AE_FULLADDER_4BIT</type>
<position>121,137.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_2</ID>220 </input>
<input>
<ID>IN_3</ID>217 </input>
<output>
<ID>OUT_0</ID>231 </output>
<output>
<ID>OUT_1</ID>228 </output>
<output>
<ID>OUT_2</ID>229 </output>
<output>
<ID>OUT_3</ID>230 </output>
<input>
<ID>carry_in</ID>221 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>116,114.5</position>
<gparam>LABEL_TEXT PCOut</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>DE_TO</type>
<position>41,40</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRsend</lparam></gate>
<gate>
<ID>183</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-70,31.5</position>
<input>
<ID>ENABLE_0</ID>283 </input>
<input>
<ID>IN_0</ID>291 </input>
<input>
<ID>IN_1</ID>290 </input>
<input>
<ID>IN_2</ID>340 </input>
<input>
<ID>IN_3</ID>341 </input>
<input>
<ID>IN_4</ID>338 </input>
<input>
<ID>IN_5</ID>337 </input>
<input>
<ID>IN_6</ID>336 </input>
<input>
<ID>IN_7</ID>284 </input>
<output>
<ID>OUT_0</ID>232 </output>
<output>
<ID>OUT_1</ID>233 </output>
<output>
<ID>OUT_2</ID>234 </output>
<output>
<ID>OUT_3</ID>235 </output>
<output>
<ID>OUT_4</ID>278 </output>
<output>
<ID>OUT_5</ID>279 </output>
<output>
<ID>OUT_6</ID>280 </output>
<output>
<ID>OUT_7</ID>281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>-121,58</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>-120.5,29</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>-34.5,70.5</position>
<gparam>LABEL_TEXT Write MDR input into RAM at MAR address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>-31,64.5</position>
<gparam>LABEL_TEXT Write contents of RAM at MAR address to MDR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AE_REGISTER8</type>
<position>285,55</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>323 </input>
<input>
<ID>IN_2</ID>322 </input>
<input>
<ID>IN_3</ID>321 </input>
<input>
<ID>IN_4</ID>320 </input>
<input>
<ID>IN_5</ID>319 </input>
<input>
<ID>IN_6</ID>289 </input>
<input>
<ID>IN_7</ID>333 </input>
<output>
<ID>OUT_0</ID>433 </output>
<output>
<ID>OUT_1</ID>439 </output>
<output>
<ID>OUT_2</ID>147 </output>
<output>
<ID>OUT_3</ID>143 </output>
<output>
<ID>OUT_4</ID>139 </output>
<output>
<ID>OUT_5</ID>135 </output>
<output>
<ID>OUT_6</ID>339 </output>
<output>
<ID>OUT_7</ID>152 </output>
<input>
<ID>clock</ID>335 </input>
<input>
<ID>load</ID>160 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>214</ID>
<type>AE_REGISTER8</type>
<position>-61.5,129.5</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>304 </input>
<input>
<ID>IN_2</ID>305 </input>
<input>
<ID>IN_3</ID>306 </input>
<input>
<ID>IN_4</ID>307 </input>
<input>
<ID>IN_5</ID>308 </input>
<input>
<ID>IN_6</ID>309 </input>
<input>
<ID>IN_7</ID>310 </input>
<output>
<ID>OUT_0</ID>318 </output>
<output>
<ID>OUT_1</ID>317 </output>
<output>
<ID>OUT_2</ID>316 </output>
<output>
<ID>OUT_3</ID>315 </output>
<output>
<ID>OUT_4</ID>314 </output>
<output>
<ID>OUT_5</ID>313 </output>
<output>
<ID>OUT_6</ID>312 </output>
<output>
<ID>OUT_7</ID>311 </output>
<input>
<ID>clear</ID>302 </input>
<input>
<ID>clock</ID>335 </input>
<input>
<ID>load</ID>301 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>-69.5,151</position>
<gparam>LABEL_TEXT Global Bus</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_TOGGLE</type>
<position>-62.5,139.5</position>
<output>
<ID>OUT_0</ID>301 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>-63,143</position>
<gparam>LABEL_TEXT Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_TOGGLE</type>
<position>-60.5,121</position>
<output>
<ID>OUT_0</ID>302 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>-60,118.5</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_LABEL</type>
<position>218.5,121</position>
<gparam>LABEL_TEXT SR2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>-81.5,138.5</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 7</lparam></gate>
<gate>
<ID>225</ID>
<type>DA_FROM</type>
<position>-81,135</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 6</lparam></gate>
<gate>
<ID>226</ID>
<type>DA_FROM</type>
<position>-81.5,131.5</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 5</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>-81.5,128.5</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 4</lparam></gate>
<gate>
<ID>228</ID>
<type>DA_FROM</type>
<position>-81.5,125</position>
<input>
<ID>IN_0</ID>306 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 3</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>-81.5,121.5</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 2</lparam></gate>
<gate>
<ID>230</ID>
<type>DA_FROM</type>
<position>-81.5,118</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 1</lparam></gate>
<gate>
<ID>231</ID>
<type>DA_FROM</type>
<position>-81.5,114.5</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 0</lparam></gate>
<gate>
<ID>232</ID>
<type>AE_REGISTER8</type>
<position>286.5,31</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>323 </input>
<input>
<ID>IN_2</ID>322 </input>
<input>
<ID>IN_3</ID>321 </input>
<input>
<ID>IN_4</ID>320 </input>
<input>
<ID>IN_5</ID>319 </input>
<input>
<ID>IN_6</ID>289 </input>
<input>
<ID>IN_7</ID>333 </input>
<output>
<ID>OUT_0</ID>432 </output>
<output>
<ID>OUT_1</ID>438 </output>
<output>
<ID>OUT_2</ID>148 </output>
<output>
<ID>OUT_3</ID>144 </output>
<output>
<ID>OUT_4</ID>140 </output>
<output>
<ID>OUT_5</ID>136 </output>
<output>
<ID>OUT_6</ID>351 </output>
<output>
<ID>OUT_7</ID>153 </output>
<input>
<ID>clock</ID>335 </input>
<input>
<ID>load</ID>174 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>233</ID>
<type>DE_TO</type>
<position>-47,140</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 7</lparam></gate>
<gate>
<ID>234</ID>
<type>DE_TO</type>
<position>-47,137.5</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 6</lparam></gate>
<gate>
<ID>235</ID>
<type>DE_TO</type>
<position>-47,135</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>236</ID>
<type>DE_TO</type>
<position>-47,132</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>237</ID>
<type>DE_TO</type>
<position>-47,129.5</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>238</ID>
<type>DE_TO</type>
<position>-47,126</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>239</ID>
<type>DE_TO</type>
<position>-47,123</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>240</ID>
<type>DE_TO</type>
<position>-47,120</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_MUX_4x1</type>
<position>352,81</position>
<input>
<ID>IN_0</ID>359 </input>
<input>
<ID>IN_1</ID>352 </input>
<input>
<ID>IN_2</ID>351 </input>
<input>
<ID>IN_3</ID>339 </input>
<output>
<ID>OUT</ID>360 </output>
<input>
<ID>SEL_0</ID>287 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>242</ID>
<type>AE_REGISTER8</type>
<position>286,6</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>323 </input>
<input>
<ID>IN_2</ID>322 </input>
<input>
<ID>IN_3</ID>321 </input>
<input>
<ID>IN_4</ID>320 </input>
<input>
<ID>IN_5</ID>319 </input>
<input>
<ID>IN_6</ID>289 </input>
<input>
<ID>IN_7</ID>333 </input>
<output>
<ID>OUT_0</ID>363 </output>
<output>
<ID>OUT_1</ID>437 </output>
<output>
<ID>OUT_2</ID>149 </output>
<output>
<ID>OUT_3</ID>145 </output>
<output>
<ID>OUT_4</ID>141 </output>
<output>
<ID>OUT_5</ID>137 </output>
<output>
<ID>OUT_6</ID>352 </output>
<output>
<ID>OUT_7</ID>154 </output>
<input>
<ID>clock</ID>335 </input>
<input>
<ID>load</ID>223 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>243</ID>
<type>AE_MUX_4x1</type>
<position>358,70</position>
<input>
<ID>IN_0</ID>359 </input>
<input>
<ID>IN_1</ID>352 </input>
<input>
<ID>IN_2</ID>351 </input>
<input>
<ID>IN_3</ID>339 </input>
<output>
<ID>OUT</ID>361 </output>
<input>
<ID>SEL_0</ID>155 </input>
<input>
<ID>SEL_1</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>244</ID>
<type>AE_REGISTER8</type>
<position>286,-19</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>323 </input>
<input>
<ID>IN_2</ID>322 </input>
<input>
<ID>IN_3</ID>321 </input>
<input>
<ID>IN_4</ID>320 </input>
<input>
<ID>IN_5</ID>319 </input>
<input>
<ID>IN_6</ID>289 </input>
<input>
<ID>IN_7</ID>333 </input>
<output>
<ID>OUT_0</ID>362 </output>
<output>
<ID>OUT_1</ID>436 </output>
<output>
<ID>OUT_2</ID>150 </output>
<output>
<ID>OUT_3</ID>146 </output>
<output>
<ID>OUT_4</ID>142 </output>
<output>
<ID>OUT_5</ID>138 </output>
<output>
<ID>OUT_6</ID>359 </output>
<output>
<ID>OUT_7</ID>354 </output>
<input>
<ID>clock</ID>335 </input>
<input>
<ID>load</ID>285 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_LABEL</type>
<position>208.5,66</position>
<gparam>LABEL_TEXT Input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>AA_LABEL</type>
<position>192,-3.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>AA_LABEL</type>
<position>219,109.5</position>
<gparam>LABEL_TEXT SR1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>-2.5,141.5</position>
<input>
<ID>IN_0</ID>325 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 7</lparam></gate>
<gate>
<ID>250</ID>
<type>DA_FROM</type>
<position>-2,138</position>
<input>
<ID>IN_0</ID>326 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 6</lparam></gate>
<gate>
<ID>251</ID>
<type>DA_FROM</type>
<position>-2.5,134.5</position>
<input>
<ID>IN_0</ID>327 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>252</ID>
<type>DA_FROM</type>
<position>-2.5,131.5</position>
<input>
<ID>IN_0</ID>328 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>253</ID>
<type>DA_FROM</type>
<position>-2.5,128</position>
<input>
<ID>IN_0</ID>329 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>254</ID>
<type>DA_FROM</type>
<position>-2.5,124.5</position>
<input>
<ID>IN_0</ID>330 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>255</ID>
<type>DA_FROM</type>
<position>-2.5,121</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>-2.5,117.5</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>258</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>465.5,51.5</position>
<input>
<ID>IN_0</ID>434 </input>
<input>
<ID>IN_1</ID>440 </input>
<input>
<ID>IN_2</ID>133 </input>
<input>
<ID>IN_3</ID>131 </input>
<input>
<ID>IN_4</ID>129 </input>
<input>
<ID>IN_5</ID>127 </input>
<input>
<ID>IN_6</ID>360 </input>
<input>
<ID>IN_7</ID>288 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>262</ID>
<type>AE_MUX_4x1</type>
<position>418.5,-44</position>
<input>
<ID>IN_0</ID>362 </input>
<input>
<ID>IN_1</ID>363 </input>
<input>
<ID>IN_2</ID>432 </input>
<input>
<ID>IN_3</ID>433 </input>
<output>
<ID>OUT</ID>434 </output>
<input>
<ID>SEL_0</ID>287 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>264</ID>
<type>AE_MUX_4x1</type>
<position>425.5,-53.5</position>
<input>
<ID>IN_0</ID>362 </input>
<input>
<ID>IN_1</ID>363 </input>
<input>
<ID>IN_2</ID>432 </input>
<input>
<ID>IN_3</ID>433 </input>
<output>
<ID>OUT</ID>435 </output>
<input>
<ID>SEL_0</ID>155 </input>
<input>
<ID>SEL_1</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>266</ID>
<type>AE_MUX_4x1</type>
<position>395.5,-2.5</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>149 </input>
<input>
<ID>IN_2</ID>148 </input>
<input>
<ID>IN_3</ID>147 </input>
<output>
<ID>OUT</ID>133 </output>
<input>
<ID>SEL_0</ID>287 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>268</ID>
<type>AE_MUX_4x1</type>
<position>401,-13</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>149 </input>
<input>
<ID>IN_2</ID>148 </input>
<input>
<ID>IN_3</ID>147 </input>
<output>
<ID>OUT</ID>134 </output>
<input>
<ID>SEL_0</ID>155 </input>
<input>
<ID>SEL_1</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_MUX_4x1</type>
<position>406.5,-23.5</position>
<input>
<ID>IN_0</ID>436 </input>
<input>
<ID>IN_1</ID>437 </input>
<input>
<ID>IN_2</ID>438 </input>
<input>
<ID>IN_3</ID>439 </input>
<output>
<ID>OUT</ID>441 </output>
<input>
<ID>SEL_0</ID>155 </input>
<input>
<ID>SEL_1</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>272</ID>
<type>AE_MUX_4x1</type>
<position>412,-33.5</position>
<input>
<ID>IN_0</ID>436 </input>
<input>
<ID>IN_1</ID>437 </input>
<input>
<ID>IN_2</ID>438 </input>
<input>
<ID>IN_3</ID>439 </input>
<output>
<ID>OUT</ID>440 </output>
<input>
<ID>SEL_0</ID>287 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>273</ID>
<type>DE_TO</type>
<position>-12.5,48.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 7</lparam></gate>
<gate>
<ID>274</ID>
<type>DE_TO</type>
<position>-13.5,46</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 6</lparam></gate>
<gate>
<ID>275</ID>
<type>DE_TO</type>
<position>-13.5,43.5</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 5</lparam></gate>
<gate>
<ID>281</ID>
<type>DA_FROM</type>
<position>21,141.5</position>
<input>
<ID>IN_0</ID>366 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRsend</lparam></gate>
<gate>
<ID>282</ID>
<type>DE_TO</type>
<position>41,42.5</position>
<input>
<ID>IN_0</ID>367 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRwrite</lparam></gate>
<gate>
<ID>283</ID>
<type>AA_TOGGLE</type>
<position>32,129</position>
<output>
<ID>OUT_0</ID>372 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>284</ID>
<type>DE_TO</type>
<position>39.5,127</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 7</lparam></gate>
<gate>
<ID>285</ID>
<type>DE_TO</type>
<position>38.5,124.5</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 6</lparam></gate>
<gate>
<ID>286</ID>
<type>DE_TO</type>
<position>38.5,122</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 5</lparam></gate>
<gate>
<ID>287</ID>
<type>DE_TO</type>
<position>38.5,119.5</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 4</lparam></gate>
<gate>
<ID>288</ID>
<type>DE_TO</type>
<position>38.5,116.5</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 3</lparam></gate>
<gate>
<ID>289</ID>
<type>DE_TO</type>
<position>39,113.5</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 2</lparam></gate>
<gate>
<ID>290</ID>
<type>DE_TO</type>
<position>39,110.5</position>
<input>
<ID>IN_0</ID>369 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 1</lparam></gate>
<gate>
<ID>291</ID>
<type>DE_TO</type>
<position>39,107.5</position>
<input>
<ID>IN_0</ID>368 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 0</lparam></gate>
<gate>
<ID>292</ID>
<type>DA_FROM</type>
<position>180,66</position>
<input>
<ID>IN_0</ID>376 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID REGin</lparam></gate>
<gate>
<ID>293</ID>
<type>DE_TO</type>
<position>43.5,45.5</position>
<input>
<ID>IN_0</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID REGin</lparam></gate>
<gate>
<ID>296</ID>
<type>DD_KEYPAD_HEX</type>
<position>81.5,-68.5</position>
<output>
<ID>OUT_0</ID>391 </output>
<output>
<ID>OUT_1</ID>390 </output>
<output>
<ID>OUT_2</ID>389 </output>
<output>
<ID>OUT_3</ID>388 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>297</ID>
<type>DD_KEYPAD_HEX</type>
<position>81.5,-83.5</position>
<output>
<ID>OUT_0</ID>387 </output>
<output>
<ID>OUT_1</ID>386 </output>
<output>
<ID>OUT_2</ID>385 </output>
<output>
<ID>OUT_3</ID>384 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>298</ID>
<type>DD_KEYPAD_HEX</type>
<position>81.5,-98</position>
<output>
<ID>OUT_0</ID>395 </output>
<output>
<ID>OUT_1</ID>394 </output>
<output>
<ID>OUT_2</ID>393 </output>
<output>
<ID>OUT_3</ID>392 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_AND2</type>
<position>120.5,-85.5</position>
<input>
<ID>IN_0</ID>380 </input>
<input>
<ID>IN_1</ID>384 </input>
<output>
<ID>OUT</ID>404 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_AND2</type>
<position>120.5,-91</position>
<input>
<ID>IN_0</ID>381 </input>
<input>
<ID>IN_1</ID>385 </input>
<output>
<ID>OUT</ID>405 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>AA_AND2</type>
<position>120.5,-96.5</position>
<input>
<ID>IN_0</ID>382 </input>
<input>
<ID>IN_1</ID>386 </input>
<output>
<ID>OUT</ID>406 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>AA_AND2</type>
<position>120.5,-102</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>387 </input>
<output>
<ID>OUT</ID>407 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_AND2</type>
<position>120.5,-107.5</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>392 </input>
<output>
<ID>OUT</ID>408 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_AND2</type>
<position>120.5,-113</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>393 </input>
<output>
<ID>OUT</ID>409 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_AND2</type>
<position>120.5,-118</position>
<input>
<ID>IN_0</ID>390 </input>
<input>
<ID>IN_1</ID>394 </input>
<output>
<ID>OUT</ID>410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>AA_AND2</type>
<position>120.5,-123.5</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>395 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>AA_MUX_2x1</type>
<position>148,-66.5</position>
<input>
<ID>IN_0</ID>403 </input>
<input>
<ID>IN_1</ID>411 </input>
<output>
<ID>OUT</ID>413 </output>
<input>
<ID>SEL_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>308</ID>
<type>AA_MUX_2x1</type>
<position>148,-72</position>
<input>
<ID>IN_0</ID>402 </input>
<input>
<ID>IN_1</ID>410 </input>
<output>
<ID>OUT</ID>414 </output>
<input>
<ID>SEL_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_MUX_2x1</type>
<position>148,-77.5</position>
<input>
<ID>IN_0</ID>401 </input>
<input>
<ID>IN_1</ID>409 </input>
<output>
<ID>OUT</ID>415 </output>
<input>
<ID>SEL_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>310</ID>
<type>AA_MUX_2x1</type>
<position>148,-82.5</position>
<input>
<ID>IN_0</ID>400 </input>
<input>
<ID>IN_1</ID>408 </input>
<output>
<ID>OUT</ID>416 </output>
<input>
<ID>SEL_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>311</ID>
<type>AA_MUX_2x1</type>
<position>148,-93</position>
<input>
<ID>IN_0</ID>399 </input>
<input>
<ID>IN_1</ID>407 </input>
<output>
<ID>OUT</ID>417 </output>
<input>
<ID>SEL_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_MUX_2x1</type>
<position>148,-98</position>
<input>
<ID>IN_0</ID>398 </input>
<input>
<ID>IN_1</ID>406 </input>
<output>
<ID>OUT</ID>418 </output>
<input>
<ID>SEL_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>313</ID>
<type>AA_MUX_2x1</type>
<position>148,-103</position>
<input>
<ID>IN_0</ID>397 </input>
<input>
<ID>IN_1</ID>405 </input>
<output>
<ID>OUT</ID>419 </output>
<input>
<ID>SEL_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>AA_MUX_2x1</type>
<position>148,-108</position>
<input>
<ID>IN_0</ID>396 </input>
<input>
<ID>IN_1</ID>404 </input>
<output>
<ID>OUT</ID>420 </output>
<input>
<ID>SEL_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>AA_TOGGLE</type>
<position>151.5,-53</position>
<output>
<ID>OUT_0</ID>412 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>316</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>178.5,-88</position>
<input>
<ID>IN_0</ID>420 </input>
<input>
<ID>IN_1</ID>419 </input>
<input>
<ID>IN_2</ID>418 </input>
<input>
<ID>IN_3</ID>417 </input>
<input>
<ID>IN_4</ID>416 </input>
<input>
<ID>IN_5</ID>415 </input>
<input>
<ID>IN_6</ID>414 </input>
<input>
<ID>IN_7</ID>413 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 136</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>317</ID>
<type>AA_LABEL</type>
<position>71,-61.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>AA_LABEL</type>
<position>72,-90</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>319</ID>
<type>AA_LABEL</type>
<position>164.5,-52.5</position>
<gparam>LABEL_TEXT Control Signal</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>320</ID>
<type>AE_FULLADDER_4BIT</type>
<position>121,-59</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>390 </input>
<input>
<ID>IN_2</ID>389 </input>
<input>
<ID>IN_3</ID>388 </input>
<input>
<ID>IN_B_0</ID>395 </input>
<input>
<ID>IN_B_1</ID>394 </input>
<input>
<ID>IN_B_2</ID>393 </input>
<input>
<ID>IN_B_3</ID>392 </input>
<output>
<ID>OUT_0</ID>396 </output>
<output>
<ID>OUT_1</ID>397 </output>
<output>
<ID>OUT_2</ID>398 </output>
<output>
<ID>OUT_3</ID>399 </output>
<output>
<ID>carry_out</ID>379 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>321</ID>
<type>AE_FULLADDER_4BIT</type>
<position>121,-75</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>382 </input>
<input>
<ID>IN_2</ID>381 </input>
<input>
<ID>IN_3</ID>380 </input>
<input>
<ID>IN_B_0</ID>387 </input>
<input>
<ID>IN_B_1</ID>386 </input>
<input>
<ID>IN_B_2</ID>385 </input>
<input>
<ID>IN_B_3</ID>384 </input>
<output>
<ID>OUT_0</ID>400 </output>
<output>
<ID>OUT_1</ID>401 </output>
<output>
<ID>OUT_2</ID>402 </output>
<output>
<ID>OUT_3</ID>403 </output>
<input>
<ID>carry_in</ID>379 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>322</ID>
<type>DD_KEYPAD_HEX</type>
<position>81.5,-55</position>
<output>
<ID>OUT_0</ID>383 </output>
<output>
<ID>OUT_1</ID>382 </output>
<output>
<ID>OUT_2</ID>381 </output>
<output>
<ID>OUT_3</ID>380 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>338</ID>
<type>DE_TO</type>
<position>-13.5,41</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 4</lparam></gate>
<gate>
<ID>339</ID>
<type>DE_TO</type>
<position>-13.5,38</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 3</lparam></gate>
<gate>
<ID>340</ID>
<type>DE_TO</type>
<position>-13,35</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 2</lparam></gate>
<gate>
<ID>341</ID>
<type>DE_TO</type>
<position>-13,32</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 1</lparam></gate>
<gate>
<ID>342</ID>
<type>DE_TO</type>
<position>-13,29</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 0</lparam></gate>
<gate>
<ID>343</ID>
<type>BB_CLOCK</type>
<position>-17.5,100</position>
<output>
<ID>CLK</ID>335 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>344</ID>
<type>DA_FROM</type>
<position>-99.5,42</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 7</lparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>-99.5,35</position>
<input>
<ID>IN_0</ID>337 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>346</ID>
<type>DA_FROM</type>
<position>-99.5,32</position>
<input>
<ID>IN_0</ID>338 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>-99.5,28.5</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>-99.5,25</position>
<input>
<ID>IN_0</ID>340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>349</ID>
<type>DA_FROM</type>
<position>-99.5,21.5</position>
<input>
<ID>IN_0</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>350</ID>
<type>DA_FROM</type>
<position>-99.5,18</position>
<input>
<ID>IN_0</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>351</ID>
<type>DA_FROM</type>
<position>-100,38</position>
<input>
<ID>IN_0</ID>336 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 6</lparam></gate>
<gate>
<ID>352</ID>
<type>DE_TO</type>
<position>148,117.5</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 7</lparam></gate>
<gate>
<ID>353</ID>
<type>DE_TO</type>
<position>147,115</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 6</lparam></gate>
<gate>
<ID>354</ID>
<type>DE_TO</type>
<position>147,112.5</position>
<input>
<ID>IN_0</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 5</lparam></gate>
<gate>
<ID>355</ID>
<type>DE_TO</type>
<position>147,110</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 4</lparam></gate>
<gate>
<ID>356</ID>
<type>DE_TO</type>
<position>147,107</position>
<input>
<ID>IN_0</ID>346 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 3</lparam></gate>
<gate>
<ID>357</ID>
<type>DE_TO</type>
<position>147.5,104</position>
<input>
<ID>IN_0</ID>345 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 2</lparam></gate>
<gate>
<ID>358</ID>
<type>DE_TO</type>
<position>147.5,101</position>
<input>
<ID>IN_0</ID>343 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 1</lparam></gate>
<gate>
<ID>359</ID>
<type>DE_TO</type>
<position>147.5,98</position>
<input>
<ID>IN_0</ID>342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus In 0</lparam></gate>
<gate>
<ID>360</ID>
<type>AE_MUX_4x1</type>
<position>364,60</position>
<input>
<ID>IN_0</ID>138 </input>
<input>
<ID>IN_1</ID>137 </input>
<input>
<ID>IN_2</ID>136 </input>
<input>
<ID>IN_3</ID>135 </input>
<output>
<ID>OUT</ID>127 </output>
<input>
<ID>SEL_0</ID>287 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>362</ID>
<type>AA_LABEL</type>
<position>155,125</position>
<gparam>LABEL_TEXT Send PC to Bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>AE_MUX_4x1</type>
<position>369.5,49</position>
<input>
<ID>IN_0</ID>138 </input>
<input>
<ID>IN_1</ID>137 </input>
<input>
<ID>IN_2</ID>136 </input>
<input>
<ID>IN_3</ID>135 </input>
<output>
<ID>OUT</ID>128 </output>
<input>
<ID>SEL_0</ID>155 </input>
<input>
<ID>SEL_1</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>364</ID>
<type>BI_ROM_12x16</type>
<position>39,67</position>
<input>
<ID>ADDRESS_0</ID>373 </input>
<input>
<ID>ADDRESS_1</ID>374 </input>
<input>
<ID>ADDRESS_2</ID>375 </input>
<input>
<ID>ADDRESS_3</ID>353 </input>
<input>
<ID>ADDRESS_4</ID>364 </input>
<input>
<ID>ADDRESS_5</ID>365 </input>
<output>
<ID>DATA_OUT_0</ID>373 </output>
<output>
<ID>DATA_OUT_1</ID>374 </output>
<output>
<ID>DATA_OUT_10</ID>167 </output>
<output>
<ID>DATA_OUT_11</ID>442 </output>
<output>
<ID>DATA_OUT_12</ID>357 </output>
<output>
<ID>DATA_OUT_13</ID>358 </output>
<output>
<ID>DATA_OUT_14</ID>356 </output>
<output>
<ID>DATA_OUT_15</ID>355 </output>
<output>
<ID>DATA_OUT_2</ID>375 </output>
<output>
<ID>DATA_OUT_8</ID>377 </output>
<output>
<ID>DATA_OUT_9</ID>367 </output>
<input>
<ID>ENABLE_0</ID>447 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 57345</lparam>
<lparam>Address:1 49154</lparam>
<lparam>Address:2 6147</lparam>
<lparam>Address:3 25604</lparam></gate>
<gate>
<ID>365</ID>
<type>AE_MUX_4x1</type>
<position>338.5,99</position>
<input>
<ID>IN_0</ID>354 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>152 </input>
<output>
<ID>OUT</ID>288 </output>
<input>
<ID>SEL_0</ID>287 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>366</ID>
<type>AE_MUX_4x1</type>
<position>374.5,38.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>141 </input>
<input>
<ID>IN_2</ID>140 </input>
<input>
<ID>IN_3</ID>139 </input>
<output>
<ID>OUT</ID>129 </output>
<input>
<ID>SEL_0</ID>287 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>367</ID>
<type>AA_LABEL</type>
<position>197,-18.5</position>
<gparam>LABEL_TEXT DR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>368</ID>
<type>AE_MUX_4x1</type>
<position>380,28.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>141 </input>
<input>
<ID>IN_2</ID>140 </input>
<input>
<ID>IN_3</ID>139 </input>
<output>
<ID>OUT</ID>130 </output>
<input>
<ID>SEL_0</ID>155 </input>
<input>
<ID>SEL_1</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>369</ID>
<type>AE_MUX_4x1</type>
<position>385.5,18</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>144 </input>
<input>
<ID>IN_3</ID>143 </input>
<output>
<ID>OUT</ID>131 </output>
<input>
<ID>SEL_0</ID>287 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>370</ID>
<type>AE_MUX_4x1</type>
<position>391,7.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>144 </input>
<input>
<ID>IN_3</ID>143 </input>
<output>
<ID>OUT</ID>132 </output>
<input>
<ID>SEL_0</ID>155 </input>
<input>
<ID>SEL_1</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>371</ID>
<type>AA_TOGGLE</type>
<position>201.5,-18</position>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>372</ID>
<type>DE_TO</type>
<position>34,21.5</position>
<input>
<ID>IN_0</ID>355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID sendPC</lparam></gate>
<gate>
<ID>374</ID>
<type>DA_FROM</type>
<position>137,128.5</position>
<input>
<ID>IN_0</ID>344 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID sendPC</lparam></gate>
<gate>
<ID>375</ID>
<type>DA_FROM</type>
<position>-99,70.5</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 7</lparam></gate>
<gate>
<ID>376</ID>
<type>DA_FROM</type>
<position>-99,63.5</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 5</lparam></gate>
<gate>
<ID>377</ID>
<type>DA_FROM</type>
<position>-99,60.5</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 4</lparam></gate>
<gate>
<ID>378</ID>
<type>DA_FROM</type>
<position>-99,57</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 3</lparam></gate>
<gate>
<ID>379</ID>
<type>DA_FROM</type>
<position>-99,53.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 2</lparam></gate>
<gate>
<ID>380</ID>
<type>DA_FROM</type>
<position>-99,50</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 1</lparam></gate>
<gate>
<ID>381</ID>
<type>DA_FROM</type>
<position>-99,46.5</position>
<input>
<ID>IN_0</ID>202 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 0</lparam></gate>
<gate>
<ID>382</ID>
<type>DA_FROM</type>
<position>-99,66.5</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus Out 6</lparam></gate>
<gate>
<ID>383</ID>
<type>BA_DECODER_2x4</type>
<position>212,-11.5</position>
<input>
<ID>ENABLE</ID>376 </input>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT_0</ID>285 </output>
<output>
<ID>OUT_1</ID>223 </output>
<output>
<ID>OUT_2</ID>174 </output>
<output>
<ID>OUT_3</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>DA_FROM</type>
<position>-61,69.5</position>
<input>
<ID>IN_0</ID>283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDRwrite</lparam></gate>
<gate>
<ID>385</ID>
<type>AE_MUX_4x1</type>
<position>344.5,89.5</position>
<input>
<ID>IN_0</ID>354 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>152 </input>
<output>
<ID>OUT</ID>334 </output>
<input>
<ID>SEL_0</ID>155 </input>
<input>
<ID>SEL_1</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>-49.5,62</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID MAR</lparam></gate>
<gate>
<ID>388</ID>
<type>DE_TO</type>
<position>34.5,25</position>
<input>
<ID>IN_0</ID>356 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR</lparam></gate>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-112,95.5,-63</points>
<intersection>-112 3</intersection>
<intersection>-67.5 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-63,117,-63</points>
<connection>
<GID>320</GID>
<name>IN_2</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-67.5,95.5,-67.5</points>
<connection>
<GID>296</GID>
<name>OUT_2</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>95.5,-112,117.5,-112</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-117,94.5,-62</points>
<intersection>-117 3</intersection>
<intersection>-69.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94.5,-62,117,-62</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>94.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-69.5,94.5,-69.5</points>
<connection>
<GID>296</GID>
<name>OUT_1</name></connection>
<intersection>94.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>94.5,-117,117.5,-117</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-107.5,-27.5,-106.5,-27.5</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-106.5,-27.5,-106.5,-26</points>
<intersection>-27.5 1</intersection>
<intersection>-26 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-106.5,-26,-105.5,-26</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-106.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-122.5,93.5,-61</points>
<intersection>-122.5 3</intersection>
<intersection>-71.5 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-61,117,-61</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-71.5,93.5,-71.5</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>93.5,-122.5,117.5,-122.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-29.5,-106.5,-29</points>
<intersection>-29.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-106.5,-29,-105.5,-29</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-107.5,-29.5,-106.5,-29.5</points>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-108.5,103,-57</points>
<intersection>-108.5 3</intersection>
<intersection>-95 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-57,117,-57</points>
<connection>
<GID>320</GID>
<name>IN_B_3</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-95,103,-95</points>
<connection>
<GID>298</GID>
<name>OUT_3</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103,-108.5,117.5,-108.5</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106.5,-32,-106.5,-31.5</points>
<intersection>-32 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-106.5,-32,-105.5,-32</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-107.5,-31.5,-106.5,-31.5</points>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>-106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-114,102.5,-56</points>
<intersection>-114 3</intersection>
<intersection>-97 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-56,117,-56</points>
<connection>
<GID>320</GID>
<name>IN_B_2</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-97,102.5,-97</points>
<connection>
<GID>298</GID>
<name>OUT_2</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,-114,117.5,-114</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-107.5,-33.5,-106.5,-33.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-106.5,-47,-106.5,-33.5</points>
<intersection>-47 8</intersection>
<intersection>-44 9</intersection>
<intersection>-41 10</intersection>
<intersection>-38 11</intersection>
<intersection>-35 12</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-106.5,-47,-105.5,-47</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-106.5,-44,-105.5,-44</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-106.5,-41,-105.5,-41</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-106.5,-38,-105.5,-38</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-106.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-106.5,-35,-105.5,-35</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-106.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-119,102,-55</points>
<intersection>-119 3</intersection>
<intersection>-99 2</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-55,117,-55</points>
<connection>
<GID>320</GID>
<name>IN_B_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-99,102,-99</points>
<connection>
<GID>298</GID>
<name>OUT_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102,-119,117.5,-119</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-38.5,-59.5,-35.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-35.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-59.5,-35.5,-59,-35.5</points>
<intersection>-59.5 0</intersection>
<intersection>-59 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-59,-35.5,-59,-34.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-35.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-124.5,101,-54</points>
<intersection>-124.5 3</intersection>
<intersection>-101 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-54,117,-54</points>
<connection>
<GID>320</GID>
<name>IN_B_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-101,101,-101</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101,-124.5,117.5,-124.5</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-38.5,-60.5,-35.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-62,-35.5,-60.5,-35.5</points>
<intersection>-62 4</intersection>
<intersection>-60.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-62,-35.5,-62,-34.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-35.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-109,137,-57.5</points>
<intersection>-109 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-109,146,-109</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-57.5,137,-57.5</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-65,-36.5,-61.5,-36.5</points>
<intersection>-65 4</intersection>
<intersection>-61.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-61.5,-38.5,-61.5,-36.5</points>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<intersection>-36.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-65,-36.5,-65,-34.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-36.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-104,136,-58.5</points>
<intersection>-104 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-104,146,-104</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-58.5,136,-58.5</points>
<connection>
<GID>320</GID>
<name>OUT_1</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-68,-37.5,-62.5,-37.5</points>
<intersection>-68 5</intersection>
<intersection>-62.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-62.5,-38.5,-62.5,-37.5</points>
<connection>
<GID>15</GID>
<name>IN_3</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-68,-37.5,-68,-34.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-37.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-99,135,-59.5</points>
<intersection>-99 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-99,146,-99</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-59.5,135,-59.5</points>
<connection>
<GID>320</GID>
<name>OUT_2</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-47,-37.5,-47,-34.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-37.5,-47,-37.5</points>
<intersection>-52.5 3</intersection>
<intersection>-47 1</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-52.5,-38.5,-52.5,-37.5</points>
<connection>
<GID>15</GID>
<name>IN_B_0</name></connection>
<intersection>-37.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-94,134,-60.5</points>
<intersection>-94 1</intersection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-94,146,-94</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-60.5,134,-60.5</points>
<connection>
<GID>320</GID>
<name>OUT_3</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,-38.5,-53.5,-36.5</points>
<connection>
<GID>15</GID>
<name>IN_B_1</name></connection>
<intersection>-36.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-50,-36.5,-50,-34.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-36.5,-50,-36.5</points>
<intersection>-53.5 0</intersection>
<intersection>-50 1</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-83.5,133,-73.5</points>
<intersection>-83.5 1</intersection>
<intersection>-73.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-83.5,146,-83.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-73.5,133,-73.5</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53,-35.5,-53,-34.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-54.5,-38.5,-54.5,-35.5</points>
<connection>
<GID>15</GID>
<name>IN_B_2</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-54.5,-35.5,-53,-35.5</points>
<intersection>-54.5 1</intersection>
<intersection>-53 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-78.5,132,-74.5</points>
<intersection>-78.5 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-78.5,146,-78.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-74.5,132,-74.5</points>
<connection>
<GID>321</GID>
<name>OUT_1</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-55.5,-38.5,-55.5,-35.5</points>
<connection>
<GID>15</GID>
<name>IN_B_3</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-56,-35.5,-55.5,-35.5</points>
<intersection>-56 4</intersection>
<intersection>-55.5 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-56,-35.5,-56,-34.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-35.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-75.5,131,-73</points>
<intersection>-75.5 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,-73,146,-73</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-75.5,131,-75.5</points>
<connection>
<GID>321</GID>
<name>OUT_2</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-38.5,-1.5,-35.5</points>
<connection>
<GID>14</GID>
<name>IN_B_3</name></connection>
<intersection>-35.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2,-35.5,-1.5,-35.5</points>
<intersection>-2 5</intersection>
<intersection>-1.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-2,-35.5,-2,-34.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-35.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-76.5,130,-67.5</points>
<intersection>-76.5 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-67.5,146,-67.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-76.5,130,-76.5</points>
<connection>
<GID>321</GID>
<name>OUT_3</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-35.5,1,-34.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-0.5,-38.5,-0.5,-35.5</points>
<connection>
<GID>14</GID>
<name>IN_B_2</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-35.5,1,-35.5</points>
<intersection>-0.5 1</intersection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-107,132.5,-85.5</points>
<intersection>-107 1</intersection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-107,146,-107</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-85.5,132.5,-85.5</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-38.5,0.5,-36.5</points>
<connection>
<GID>14</GID>
<name>IN_B_1</name></connection>
<intersection>-36.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>4,-36.5,4,-34.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>0.5,-36.5,4,-36.5</points>
<intersection>0.5 0</intersection>
<intersection>4 1</intersection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-102,131.5,-91</points>
<intersection>-102 1</intersection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-102,146,-102</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>131.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-91,131.5,-91</points>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-38.5,1.5,-37.5</points>
<connection>
<GID>14</GID>
<name>IN_B_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>7,-37.5,7,-34.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-37.5,7,-37.5</points>
<intersection>1.5 0</intersection>
<intersection>7 1</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-97,130.5,-96.5</points>
<intersection>-97 1</intersection>
<intersection>-96.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-97,146,-97</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-96.5,130.5,-96.5</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-38.5,-5.5,-35.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-5,-35.5,-5,-34.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,-35.5,-5,-35.5</points>
<intersection>-5.5 0</intersection>
<intersection>-5 1</intersection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-102,130.5,-92</points>
<intersection>-102 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-92,146,-92</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-102,130.5,-102</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,-38.5,-6.5,-35.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-8,-35.5,-8,-34.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8,-35.5,-6.5,-35.5</points>
<intersection>-8 1</intersection>
<intersection>-6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-107.5,129.5,-81.5</points>
<intersection>-107.5 2</intersection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-81.5,146,-81.5</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-107.5,129.5,-107.5</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-38.5,-7.5,-36.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>-36.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-11,-36.5,-11,-34.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-11,-36.5,-7.5,-36.5</points>
<intersection>-11 1</intersection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-113.5,134,-76.5</points>
<intersection>-113.5 2</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-76.5,146,-76.5</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-113.5,134,-113.5</points>
<intersection>123.5 3</intersection>
<intersection>134 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>123.5,-113.5,123.5,-113</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<intersection>-113.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-14,-37.5,-14,-34.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14,-37.5,-8.5,-37.5</points>
<intersection>-14 1</intersection>
<intersection>-8.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-8.5,-38.5,-8.5,-37.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>-37.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-118,134.5,-71</points>
<intersection>-118 2</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134.5,-71,146,-71</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>134.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-118,134.5,-118</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<intersection>134.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>-10,-48.5,-4,-48.5</points>
<intersection>-10 13</intersection>
<intersection>-4 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-4,-48.5,-4,-46.5</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<intersection>-48.5 11</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-10,-56.5,-10,-48.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>-48.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-123.5,135,-65.5</points>
<intersection>-123.5 2</intersection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-65.5,146,-65.5</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-123.5,135,-123.5</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-53.5,3,-48.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>-48.5 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-3,-48.5,3,-48.5</points>
<intersection>-3 17</intersection>
<intersection>3 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>-3,-48.5,-3,-46.5</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<intersection>-48.5 16</intersection></vsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-105.5,148,-53</points>
<connection>
<GID>314</GID>
<name>SEL_0</name></connection>
<connection>
<GID>313</GID>
<name>SEL_0</name></connection>
<connection>
<GID>312</GID>
<name>SEL_0</name></connection>
<connection>
<GID>311</GID>
<name>SEL_0</name></connection>
<connection>
<GID>310</GID>
<name>SEL_0</name></connection>
<connection>
<GID>309</GID>
<name>SEL_0</name></connection>
<connection>
<GID>308</GID>
<name>SEL_0</name></connection>
<connection>
<GID>307</GID>
<name>SEL_0</name></connection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148,-53,149.5,-53</points>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-47.5,-2,-46.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-2,-47.5,17,-47.5</points>
<intersection>-2 0</intersection>
<intersection>17 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17,-50.5,17,-47.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>-47.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-84,173.5,-66.5</points>
<connection>
<GID>316</GID>
<name>IN_7</name></connection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>150,-66.5,173.5,-66.5</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-49.5,15,-49.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>15 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>15,-50.5,15,-49.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-49.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-85,172,-72</points>
<intersection>-85 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172,-85,173.5,-85</points>
<connection>
<GID>316</GID>
<name>IN_6</name></connection>
<intersection>172 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150,-72,172,-72</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76,-73.5,19.5,-73.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 34</intersection>
<intersection>-50 32</intersection>
<intersection>-37 28</intersection>
<intersection>-23 22</intersection>
<intersection>-9.5 13</intersection>
<intersection>3.5 8</intersection>
<intersection>17.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>17.5,-73.5,17.5,-52.5</points>
<intersection>-73.5 1</intersection>
<intersection>-52.5 38</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>3.5,-73.5,3.5,-55.5</points>
<intersection>-73.5 1</intersection>
<intersection>-55.5 42</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-9.5,-73.5,-9.5,-58.5</points>
<intersection>-73.5 1</intersection>
<intersection>-58.5 36</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>-23,-73.5,-23,-61.5</points>
<intersection>-73.5 1</intersection>
<intersection>-61.5 40</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>-37,-73.5,-37,-64.5</points>
<intersection>-73.5 1</intersection>
<intersection>-64.5 44</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>-50,-73.5,-50,-67.5</points>
<intersection>-73.5 1</intersection>
<intersection>-67.5 37</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>-63.5,-73.5,-63.5,-70.5</points>
<intersection>-73.5 1</intersection>
<intersection>-70.5 41</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>-9.5,-58.5,-8.5,-58.5</points>
<connection>
<GID>16</GID>
<name>SEL_0</name></connection>
<intersection>-9.5 13</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-50,-67.5,-49,-67.5</points>
<connection>
<GID>18</GID>
<name>SEL_0</name></connection>
<intersection>-50 32</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>17.5,-52.5,18.5,-52.5</points>
<connection>
<GID>19</GID>
<name>SEL_0</name></connection>
<intersection>17.5 4</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>-23,-61.5,-22,-61.5</points>
<connection>
<GID>21</GID>
<name>SEL_0</name></connection>
<intersection>-23 22</intersection></hsegment>
<hsegment>
<ID>41</ID>
<points>-63.5,-70.5,-62.5,-70.5</points>
<connection>
<GID>22</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 34</intersection></hsegment>
<hsegment>
<ID>42</ID>
<points>3.5,-55.5,4.5,-55.5</points>
<connection>
<GID>23</GID>
<name>SEL_0</name></connection>
<intersection>3.5 8</intersection></hsegment>
<hsegment>
<ID>44</ID>
<points>-37,-64.5,-35.5,-64.5</points>
<connection>
<GID>17</GID>
<name>SEL_0</name></connection>
<intersection>-37 28</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-86,170.5,-77.5</points>
<intersection>-86 1</intersection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170.5,-86,173.5,-86</points>
<connection>
<GID>316</GID>
<name>IN_5</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150,-77.5,170.5,-77.5</points>
<connection>
<GID>309</GID>
<name>OUT</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-76.5,16,-54.5</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-87,169.5,-82.5</points>
<intersection>-87 1</intersection>
<intersection>-82.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-87,173.5,-87</points>
<connection>
<GID>316</GID>
<name>IN_4</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150,-82.5,169.5,-82.5</points>
<connection>
<GID>310</GID>
<name>OUT</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-53.5,1,-50.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>0.5,-50.5,1,-50.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-93,169.5,-88</points>
<intersection>-93 2</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-88,173.5,-88</points>
<connection>
<GID>316</GID>
<name>IN_3</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150,-93,169.5,-93</points>
<connection>
<GID>311</GID>
<name>OUT</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-76.5,2,-57.5</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-98,170.5,-89</points>
<intersection>-98 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170.5,-89,173.5,-89</points>
<connection>
<GID>316</GID>
<name>IN_2</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150,-98,170.5,-98</points>
<connection>
<GID>312</GID>
<name>OUT</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-59.5,-23.5,-47.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-47.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-5,-47.5,-5,-46.5</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-23.5,-47.5,-5,-47.5</points>
<intersection>-23.5 0</intersection>
<intersection>-5 1</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-103,172,-90</points>
<intersection>-103 2</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172,-90,173.5,-90</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>172 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150,-103,172,-103</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-56.5,-12,-49.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-13,-49.5,-12,-49.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-108,173.5,-91</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>150,-108,173.5,-108</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-76.5,-11,-60.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,-76.5,-24.5,-63.5</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-59.5,-25.5,-48.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-26.5,-48.5,-25.5,-48.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-62.5,-39,-49.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-40,-49.5,-39,-49.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-39 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-62.5,-37,-47.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>-47.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-56,-47.5,-56,-46.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-56,-47.5,-37,-47.5</points>
<intersection>-56 1</intersection>
<intersection>-37 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-76.5,-38,-66.5</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50.5,-65.5,-50.5,-48.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-48.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-57,-48.5,-50.5,-48.5</points>
<intersection>-57 4</intersection>
<intersection>-50.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-57,-48.5,-57,-46.5</points>
<connection>
<GID>15</GID>
<name>OUT_1</name></connection>
<intersection>-48.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-48.5,-58,-46.5</points>
<connection>
<GID>15</GID>
<name>OUT_2</name></connection>
<intersection>-48.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-64,-68.5,-64,-48.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-64,-48.5,-58,-48.5</points>
<intersection>-64 1</intersection>
<intersection>-58 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59,-47.5,-59,-46.5</points>
<connection>
<GID>15</GID>
<name>OUT_3</name></connection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-47.5,-59,-47.5</points>
<intersection>-77.5 3</intersection>
<intersection>-59 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-77.5,-71.5,-77.5,-47.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-47.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52.5,-65.5,-52.5,-50.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-50.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-53.5,-50.5,-52.5,-50.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,-68.5,-66,-49.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-49.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-67,-49.5,-66,-49.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-79.5,-71.5,-79.5,-48.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-48.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-80.5,-48.5,-79.5,-48.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329,-52.5,329,28</points>
<intersection>-52.5 2</intersection>
<intersection>28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,28,329,28</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>329 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>329,-52.5,422.5,-52.5</points>
<connection>
<GID>264</GID>
<name>IN_2</name></connection>
<intersection>329 0</intersection>
<intersection>409.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>409.5,-52.5,409.5,-43</points>
<intersection>-52.5 2</intersection>
<intersection>-43 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>409.5,-43,415.5,-43</points>
<connection>
<GID>262</GID>
<name>IN_2</name></connection>
<intersection>409.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-76.5,-51.5,-69.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,-50.5,337.5,52</points>
<intersection>-50.5 2</intersection>
<intersection>52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,52,337.5,52</points>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection>
<intersection>337.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>337.5,-50.5,422.5,-50.5</points>
<connection>
<GID>264</GID>
<name>IN_3</name></connection>
<intersection>337.5 0</intersection>
<intersection>407.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>407.5,-50.5,407.5,-41</points>
<intersection>-50.5 2</intersection>
<intersection>-41 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>407.5,-41,415.5,-41</points>
<connection>
<GID>262</GID>
<name>IN_3</name></connection>
<intersection>407.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-76.5,-65,-72.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429,-44,429,48.5</points>
<intersection>-44 2</intersection>
<intersection>48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429,48.5,460.5,48.5</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>429 0</intersection>
<intersection>460.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,-44,429,-44</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<intersection>429 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>460.5,35,460.5,48.5</points>
<intersection>35 4</intersection>
<intersection>48.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>460.5,35,479.5,35</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>460.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-78.5,-76.5,-78.5,-75.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>438.5,-53.5,438.5,8</points>
<intersection>-53.5 8</intersection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>438.5,8,462.5,8</points>
<intersection>438.5 0</intersection>
<intersection>462.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>462.5,-3.5,462.5,10.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-3.5 5</intersection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>462.5,-3.5,481.5,-3.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>462.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>428.5,-53.5,438.5,-53.5</points>
<connection>
<GID>264</GID>
<name>OUT</name></connection>
<intersection>438.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49.5,-41.5,-11.5,-41.5</points>
<connection>
<GID>14</GID>
<name>carry_out</name></connection>
<connection>
<GID>15</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,-36.5,349.5,-21</points>
<intersection>-36.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-21,349.5,-21</points>
<connection>
<GID>244</GID>
<name>OUT_1</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349.5,-36.5,409,-36.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>349.5 0</intersection>
<intersection>400.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>400.5,-36.5,400.5,-26.5</points>
<intersection>-36.5 2</intersection>
<intersection>-26.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>400.5,-26.5,403.5,-26.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>400.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,-34.5,349.5,4</points>
<intersection>-34.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,4,349.5,4</points>
<connection>
<GID>242</GID>
<name>OUT_1</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349.5,-34.5,409,-34.5</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<intersection>349.5 0</intersection>
<intersection>398 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>398,-34.5,398,-24.5</points>
<intersection>-34.5 2</intersection>
<intersection>-24.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>398,-24.5,403.5,-24.5</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<intersection>398 3</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,-32.5,349.5,29</points>
<intersection>-32.5 2</intersection>
<intersection>29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,29,349.5,29</points>
<connection>
<GID>232</GID>
<name>OUT_1</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349.5,-32.5,409,-32.5</points>
<connection>
<GID>272</GID>
<name>IN_2</name></connection>
<intersection>349.5 0</intersection>
<intersection>395.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>395.5,-32.5,395.5,-22.5</points>
<intersection>-32.5 2</intersection>
<intersection>-22.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>395.5,-22.5,403.5,-22.5</points>
<connection>
<GID>270</GID>
<name>IN_2</name></connection>
<intersection>395.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,-30.5,349.5,53</points>
<intersection>-30.5 2</intersection>
<intersection>53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,53,349.5,53</points>
<connection>
<GID>189</GID>
<name>OUT_1</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349.5,-30.5,409,-30.5</points>
<connection>
<GID>272</GID>
<name>IN_3</name></connection>
<intersection>349.5 0</intersection>
<intersection>393 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>393,-30.5,393,-20.5</points>
<intersection>-30.5 2</intersection>
<intersection>-20.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>393,-20.5,403.5,-20.5</points>
<connection>
<GID>270</GID>
<name>IN_3</name></connection>
<intersection>393 3</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437.5,-33.5,437.5,49.5</points>
<intersection>-33.5 2</intersection>
<intersection>49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>437.5,49.5,460.5,49.5</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<intersection>437.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>415,-33.5,437.5,-33.5</points>
<connection>
<GID>272</GID>
<name>OUT</name></connection>
<intersection>437.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436,-23.5,436,11.5</points>
<intersection>-23.5 2</intersection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436,11.5,462.5,11.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>436 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>409.5,-23.5,436,-23.5</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>436 0</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,37.5,35.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_11</name></connection>
<intersection>37.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>35.5,37.5,35.5,37.5</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,131.5,34,131.5</points>
<connection>
<GID>129</GID>
<name>OUT_4</name></connection>
<connection>
<GID>409</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,114,99.5,121.5</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>114 2</intersection>
<intersection>116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,116,101,116</points>
<connection>
<GID>411</GID>
<name>OUT_0</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,114,101,114</points>
<connection>
<GID>154</GID>
<name>count_enable</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,115,104,116</points>
<connection>
<GID>415</GID>
<name>OUT_0</name></connection>
<intersection>115 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>102,114,102,115</points>
<connection>
<GID>154</GID>
<name>count_up</name></connection>
<intersection>115 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>102,115,104,115</points>
<intersection>102 1</intersection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,98.5,103.5,103</points>
<intersection>98.5 2</intersection>
<intersection>103 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>108,98.5,108,99</points>
<connection>
<GID>424</GID>
<name>OUT_0</name></connection>
<intersection>98.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>103.5,98.5,108,98.5</points>
<intersection>103.5 0</intersection>
<intersection>108 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102,103,103.5,103</points>
<connection>
<GID>154</GID>
<name>clear</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,66.5,48,87</points>
<connection>
<GID>364</GID>
<name>ENABLE_0</name></connection>
<intersection>87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,87,48.5,87</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,57,-53.5,62</points>
<intersection>57 1</intersection>
<intersection>62 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,57,-53.5,57</points>
<connection>
<GID>147</GID>
<name>ENABLE_0</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-53.5,62,-51.5,62</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>-53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>185.5,20,185.5,35.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>20 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>178,20,185.5,20</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>185.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,28,184,36.5</points>
<intersection>28 2</intersection>
<intersection>36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,36.5,185.5,36.5</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,28,184,28</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,33,182.5,37.5</points>
<intersection>33 1</intersection>
<intersection>37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,33,182.5,33</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>182.5,37.5,185.5,37.5</points>
<connection>
<GID>95</GID>
<name>IN_2</name></connection>
<intersection>182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,38.5,185.5,38.5</points>
<connection>
<GID>95</GID>
<name>IN_3</name></connection>
<connection>
<GID>111</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,39.5,177,42.5</points>
<intersection>39.5 1</intersection>
<intersection>42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,39.5,185.5,39.5</points>
<connection>
<GID>95</GID>
<name>IN_4</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157,42.5,177,42.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,40.5,178.5,44.5</points>
<intersection>40.5 1</intersection>
<intersection>44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,40.5,185.5,40.5</points>
<connection>
<GID>95</GID>
<name>IN_5</name></connection>
<intersection>178.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>158,44.5,178.5,44.5</points>
<intersection>158 3</intersection>
<intersection>178.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>158,44.5,158,48</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>44.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,41.5,181.5,52</points>
<intersection>41.5 1</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181.5,41.5,185.5,41.5</points>
<connection>
<GID>95</GID>
<name>IN_6</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,52,181.5,52</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,42.5,184,56</points>
<intersection>42.5 1</intersection>
<intersection>56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,42.5,185.5,42.5</points>
<connection>
<GID>95</GID>
<name>IN_7</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,56,184,56</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-44.5,39,-44.5,39.5</points>
<connection>
<GID>118</GID>
<name>clear</name></connection>
<intersection>39 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-46.5,39,-44.5,39</points>
<intersection>-46.5 11</intersection>
<intersection>-44.5 4</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-46.5,38,-46.5,39</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>39 10</intersection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,50,-32,52.5</points>
<connection>
<GID>148</GID>
<name>ENABLE_0</name></connection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,52.5,-31,52.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>-32 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,48.5,-34,48.5</points>
<connection>
<GID>118</GID>
<name>OUT_7</name></connection>
<connection>
<GID>148</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,47.5,-34,47.5</points>
<connection>
<GID>118</GID>
<name>OUT_6</name></connection>
<connection>
<GID>148</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,46.5,-34,46.5</points>
<connection>
<GID>118</GID>
<name>OUT_5</name></connection>
<connection>
<GID>148</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,45.5,-34,45.5</points>
<connection>
<GID>118</GID>
<name>OUT_4</name></connection>
<connection>
<GID>148</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,44.5,-34,44.5</points>
<connection>
<GID>118</GID>
<name>OUT_3</name></connection>
<connection>
<GID>148</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,43.5,-34,43.5</points>
<connection>
<GID>118</GID>
<name>OUT_2</name></connection>
<connection>
<GID>148</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413.5,53.5,413.5,60</points>
<intersection>53.5 1</intersection>
<intersection>60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>413.5,53.5,460.5,53.5</points>
<connection>
<GID>258</GID>
<name>IN_5</name></connection>
<intersection>413.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>367,60,413.5,60</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<intersection>413.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>417.5,15.5,417.5,49</points>
<intersection>15.5 1</intersection>
<intersection>49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>417.5,15.5,462.5,15.5</points>
<connection>
<GID>101</GID>
<name>IN_5</name></connection>
<intersection>417.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,49,417.5,49</points>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<intersection>417.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>419,38.5,419,52.5</points>
<intersection>38.5 2</intersection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>419,52.5,460.5,52.5</points>
<connection>
<GID>258</GID>
<name>IN_4</name></connection>
<intersection>419 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>377.5,38.5,419,38.5</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<intersection>419 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422.5,14.5,422.5,28.5</points>
<intersection>14.5 1</intersection>
<intersection>28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>422.5,14.5,462.5,14.5</points>
<connection>
<GID>101</GID>
<name>IN_4</name></connection>
<intersection>422.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>383,28.5,422.5,28.5</points>
<connection>
<GID>368</GID>
<name>OUT</name></connection>
<intersection>422.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424.5,18,424.5,51.5</points>
<intersection>18 2</intersection>
<intersection>51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>424.5,51.5,460.5,51.5</points>
<connection>
<GID>258</GID>
<name>IN_3</name></connection>
<intersection>424.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>388.5,18,424.5,18</points>
<connection>
<GID>369</GID>
<name>OUT</name></connection>
<intersection>424.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428,7.5,428,13.5</points>
<intersection>7.5 2</intersection>
<intersection>13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428,13.5,462.5,13.5</points>
<connection>
<GID>101</GID>
<name>IN_3</name></connection>
<intersection>428 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>394,7.5,428,7.5</points>
<connection>
<GID>370</GID>
<name>OUT</name></connection>
<intersection>428 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,-2.5,429.5,50.5</points>
<intersection>-2.5 2</intersection>
<intersection>50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429.5,50.5,460.5,50.5</points>
<connection>
<GID>258</GID>
<name>IN_2</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>398.5,-2.5,429.5,-2.5</points>
<connection>
<GID>266</GID>
<name>OUT</name></connection>
<intersection>429.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433,-13,433,12.5</points>
<intersection>-13 2</intersection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>433,12.5,462.5,12.5</points>
<connection>
<GID>101</GID>
<name>IN_2</name></connection>
<intersection>433 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>404,-13,433,-13</points>
<connection>
<GID>268</GID>
<name>OUT</name></connection>
<intersection>433 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,57,304,63</points>
<intersection>57 1</intersection>
<intersection>63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,57,304,57</points>
<connection>
<GID>189</GID>
<name>OUT_5</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,63,361,63</points>
<connection>
<GID>360</GID>
<name>IN_3</name></connection>
<intersection>304 0</intersection>
<intersection>313 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>313,52,313,63</points>
<intersection>52 4</intersection>
<intersection>63 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>313,52,366.5,52</points>
<connection>
<GID>363</GID>
<name>IN_3</name></connection>
<intersection>313 3</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306,33,306,61</points>
<intersection>33 1</intersection>
<intersection>61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,33,306,33</points>
<connection>
<GID>232</GID>
<name>OUT_5</name></connection>
<intersection>306 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>306,61,361,61</points>
<connection>
<GID>360</GID>
<name>IN_2</name></connection>
<intersection>306 0</intersection>
<intersection>314.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>314.5,50,314.5,61</points>
<intersection>50 4</intersection>
<intersection>61 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>314.5,50,366.5,50</points>
<connection>
<GID>363</GID>
<name>IN_2</name></connection>
<intersection>314.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308.5,8,308.5,59</points>
<intersection>8 1</intersection>
<intersection>59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,8,308.5,8</points>
<connection>
<GID>242</GID>
<name>OUT_5</name></connection>
<intersection>308.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,59,361,59</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>308.5 0</intersection>
<intersection>316.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>316.5,48,316.5,59</points>
<intersection>48 4</intersection>
<intersection>59 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>316.5,48,366.5,48</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>316.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-17,311,57</points>
<intersection>-17 1</intersection>
<intersection>57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-17,311,-17</points>
<connection>
<GID>244</GID>
<name>OUT_5</name></connection>
<intersection>311 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>311,57,361,57</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>311 0</intersection>
<intersection>319 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>319,46,319,57</points>
<intersection>46 4</intersection>
<intersection>57 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319,46,366.5,46</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>319 3</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,41.5,312.5,56</points>
<intersection>41.5 2</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,56,312.5,56</points>
<connection>
<GID>189</GID>
<name>OUT_4</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>312.5,41.5,371.5,41.5</points>
<connection>
<GID>366</GID>
<name>IN_3</name></connection>
<intersection>312.5 0</intersection>
<intersection>319.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>319.5,31.5,319.5,41.5</points>
<intersection>31.5 4</intersection>
<intersection>41.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>319.5,31.5,377,31.5</points>
<connection>
<GID>368</GID>
<name>IN_3</name></connection>
<intersection>319.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,32,313,39.5</points>
<intersection>32 1</intersection>
<intersection>39.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,32,313,32</points>
<connection>
<GID>232</GID>
<name>OUT_4</name></connection>
<intersection>313 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,39.5,371.5,39.5</points>
<connection>
<GID>366</GID>
<name>IN_2</name></connection>
<intersection>313 0</intersection>
<intersection>321.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>321.5,29.5,321.5,39.5</points>
<intersection>29.5 4</intersection>
<intersection>39.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>321.5,29.5,377,29.5</points>
<connection>
<GID>368</GID>
<name>IN_2</name></connection>
<intersection>321.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315,7,315,37.5</points>
<intersection>7 1</intersection>
<intersection>37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,7,315,7</points>
<connection>
<GID>242</GID>
<name>OUT_4</name></connection>
<intersection>315 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>315,37.5,371.5,37.5</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>315 0</intersection>
<intersection>324 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>324,27.5,324,37.5</points>
<intersection>27.5 4</intersection>
<intersection>37.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>324,27.5,377,27.5</points>
<connection>
<GID>368</GID>
<name>IN_1</name></connection>
<intersection>324 3</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317.5,-18,317.5,35.5</points>
<intersection>-18 1</intersection>
<intersection>35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-18,317.5,-18</points>
<connection>
<GID>244</GID>
<name>OUT_4</name></connection>
<intersection>317.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>317.5,35.5,371.5,35.5</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>317.5 0</intersection>
<intersection>326.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>326.5,25.5,326.5,35.5</points>
<intersection>25.5 4</intersection>
<intersection>35.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>326.5,25.5,377,25.5</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>326.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330.5,21,330.5,55</points>
<intersection>21 2</intersection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,55,330.5,55</points>
<connection>
<GID>189</GID>
<name>OUT_3</name></connection>
<intersection>330.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>330.5,21,382.5,21</points>
<connection>
<GID>369</GID>
<name>IN_3</name></connection>
<intersection>330.5 0</intersection>
<intersection>339.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>339.5,10.5,339.5,21</points>
<intersection>10.5 4</intersection>
<intersection>21 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>339.5,10.5,388,10.5</points>
<connection>
<GID>370</GID>
<name>IN_3</name></connection>
<intersection>339.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,19,332,31</points>
<intersection>19 2</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,31,332,31</points>
<connection>
<GID>232</GID>
<name>OUT_3</name></connection>
<intersection>332 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>332,19,382.5,19</points>
<connection>
<GID>369</GID>
<name>IN_2</name></connection>
<intersection>332 0</intersection>
<intersection>342 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>342,8.5,342,19</points>
<intersection>8.5 4</intersection>
<intersection>19 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>342,8.5,388,8.5</points>
<connection>
<GID>370</GID>
<name>IN_2</name></connection>
<intersection>342 3</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>333,6,333,17</points>
<intersection>6 1</intersection>
<intersection>17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,6,333,6</points>
<connection>
<GID>242</GID>
<name>OUT_3</name></connection>
<intersection>333 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>333,17,382.5,17</points>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<intersection>333 0</intersection>
<intersection>344.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>344.5,6.5,344.5,17</points>
<intersection>6.5 4</intersection>
<intersection>17 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>344.5,6.5,388,6.5</points>
<connection>
<GID>370</GID>
<name>IN_1</name></connection>
<intersection>344.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335,-19,335,15</points>
<intersection>-19 1</intersection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-19,335,-19</points>
<connection>
<GID>244</GID>
<name>OUT_3</name></connection>
<intersection>335 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>335,15,382.5,15</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>335 0</intersection>
<intersection>347.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>347.5,4.5,347.5,15</points>
<intersection>4.5 4</intersection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>347.5,4.5,388,4.5</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>347.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370,0.5,370,54</points>
<intersection>0.5 2</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,54,370,54</points>
<connection>
<GID>189</GID>
<name>OUT_2</name></connection>
<intersection>370 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>370,0.5,392.5,0.5</points>
<connection>
<GID>266</GID>
<name>IN_3</name></connection>
<intersection>370 0</intersection>
<intersection>373.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>373.5,-10,373.5,0.5</points>
<intersection>-10 4</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>373.5,-10,398,-10</points>
<connection>
<GID>268</GID>
<name>IN_3</name></connection>
<intersection>373.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>367.5,-1.5,367.5,30</points>
<intersection>-1.5 2</intersection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,30,367.5,30</points>
<connection>
<GID>232</GID>
<name>OUT_2</name></connection>
<intersection>367.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>367.5,-1.5,392.5,-1.5</points>
<connection>
<GID>266</GID>
<name>IN_2</name></connection>
<intersection>367.5 0</intersection>
<intersection>375.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>375.5,-12,375.5,-1.5</points>
<intersection>-12 4</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>375.5,-12,398,-12</points>
<connection>
<GID>268</GID>
<name>IN_2</name></connection>
<intersection>375.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341,-3.5,341,5</points>
<intersection>-3.5 2</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,5,341,5</points>
<connection>
<GID>242</GID>
<name>OUT_2</name></connection>
<intersection>341 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341,-3.5,392.5,-3.5</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>341 0</intersection>
<intersection>378 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>378,-14,378,-3.5</points>
<intersection>-14 4</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>378,-14,398,-14</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>378 3</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341,-20,341,-5.5</points>
<intersection>-20 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-20,341,-20</points>
<connection>
<GID>244</GID>
<name>OUT_2</name></connection>
<intersection>341 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>341,-5.5,392.5,-5.5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>341 0</intersection>
<intersection>380 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>380,-16,380,-5.5</points>
<intersection>-16 4</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>380,-16,398,-16</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>380 3</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,59,290,102</points>
<intersection>59 6</intersection>
<intersection>102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,102,335.5,102</points>
<connection>
<GID>365</GID>
<name>IN_3</name></connection>
<intersection>290 0</intersection>
<intersection>303.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>303.5,92.5,303.5,102</points>
<intersection>92.5 5</intersection>
<intersection>102 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>303.5,92.5,341.5,92.5</points>
<connection>
<GID>385</GID>
<name>IN_3</name></connection>
<intersection>303.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>289,59,290,59</points>
<connection>
<GID>189</GID>
<name>OUT_7</name></connection>
<intersection>290 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291.5,35,291.5,100</points>
<intersection>35 2</intersection>
<intersection>100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>291.5,100,335.5,100</points>
<connection>
<GID>365</GID>
<name>IN_2</name></connection>
<intersection>291.5 0</intersection>
<intersection>301.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290.5,35,291.5,35</points>
<connection>
<GID>232</GID>
<name>OUT_7</name></connection>
<intersection>291.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>301.5,90.5,301.5,100</points>
<intersection>90.5 4</intersection>
<intersection>100 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>301.5,90.5,341.5,90.5</points>
<connection>
<GID>385</GID>
<name>IN_2</name></connection>
<intersection>301.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293.5,10,293.5,98</points>
<intersection>10 2</intersection>
<intersection>98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293.5,98,335.5,98</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<intersection>293.5 0</intersection>
<intersection>299.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290,10,293.5,10</points>
<connection>
<GID>242</GID>
<name>OUT_7</name></connection>
<intersection>293.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>299.5,88.5,299.5,98</points>
<intersection>88.5 4</intersection>
<intersection>98 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>299.5,88.5,341.5,88.5</points>
<connection>
<GID>385</GID>
<name>IN_1</name></connection>
<intersection>299.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426.5,-48.5,426.5,121</points>
<connection>
<GID>264</GID>
<name>SEL_0</name></connection>
<intersection>-7.5 11</intersection>
<intersection>53 5</intersection>
<intersection>71 3</intersection>
<intersection>121 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,121,426.5,121</points>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>402,71,426.5,71</points>
<intersection>402 6</intersection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>388.5,53,426.5,53</points>
<intersection>388.5 8</intersection>
<intersection>426.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>402,71,402,94.5</points>
<intersection>71 3</intersection>
<intersection>94.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>345.5,94.5,402,94.5</points>
<connection>
<GID>385</GID>
<name>SEL_0</name></connection>
<intersection>402 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>388.5,53,388.5,75.5</points>
<intersection>53 5</intersection>
<intersection>54 12</intersection>
<intersection>75.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>359,75.5,388.5,75.5</points>
<intersection>359 10</intersection>
<intersection>388.5 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>359,75,359,75.5</points>
<connection>
<GID>243</GID>
<name>SEL_0</name></connection>
<intersection>75.5 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>402,-7.5,426.5,-7.5</points>
<intersection>402 16</intersection>
<intersection>407.5 18</intersection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>370.5,54,392,54</points>
<connection>
<GID>363</GID>
<name>SEL_0</name></connection>
<intersection>388.5 8</intersection>
<intersection>392 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>392,12.5,392,54</points>
<connection>
<GID>370</GID>
<name>SEL_0</name></connection>
<intersection>35 15</intersection>
<intersection>54 12</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>381,35,392,35</points>
<intersection>381 17</intersection>
<intersection>392 13</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>402,-8,402,-7.5</points>
<connection>
<GID>268</GID>
<name>SEL_0</name></connection>
<intersection>-7.5 11</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>381,33.5,381,35</points>
<connection>
<GID>368</GID>
<name>SEL_0</name></connection>
<intersection>35 15</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>407.5,-18.5,407.5,-7.5</points>
<connection>
<GID>270</GID>
<name>SEL_0</name></connection>
<intersection>-7.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398.5,79.5,398.5,124.5</points>
<intersection>79.5 5</intersection>
<intersection>95.5 9</intersection>
<intersection>124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226.5,124.5,398.5,124.5</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>398.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>398.5,79.5,425.5,79.5</points>
<intersection>398.5 0</intersection>
<intersection>425.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>425.5,-48.5,425.5,79.5</points>
<connection>
<GID>264</GID>
<name>SEL_1</name></connection>
<intersection>-6 13</intersection>
<intersection>50 8</intersection>
<intersection>79.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>385,50,425.5,50</points>
<intersection>385 10</intersection>
<intersection>391 18</intersection>
<intersection>425.5 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>344.5,95.5,398.5,95.5</points>
<intersection>344.5 15</intersection>
<intersection>398.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>385,50,385,77</points>
<intersection>50 8</intersection>
<intersection>55.5 16</intersection>
<intersection>77 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>358,77,385,77</points>
<intersection>358 12</intersection>
<intersection>385 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>358,75,358,77</points>
<connection>
<GID>243</GID>
<name>SEL_1</name></connection>
<intersection>77 11</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>401,-6,425.5,-6</points>
<intersection>401 21</intersection>
<intersection>406.5 14</intersection>
<intersection>425.5 6</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>406.5,-18.5,406.5,-6</points>
<connection>
<GID>270</GID>
<name>SEL_1</name></connection>
<intersection>-6 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>344.5,94.5,344.5,95.5</points>
<connection>
<GID>385</GID>
<name>SEL_1</name></connection>
<intersection>95.5 9</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>369.5,55.5,385,55.5</points>
<intersection>369.5 17</intersection>
<intersection>385 10</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>369.5,54,369.5,55.5</points>
<connection>
<GID>363</GID>
<name>SEL_1</name></connection>
<intersection>55.5 16</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>391,12.5,391,50</points>
<connection>
<GID>370</GID>
<name>SEL_1</name></connection>
<intersection>36 20</intersection>
<intersection>50 8</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>380,36,391,36</points>
<intersection>380 22</intersection>
<intersection>391 18</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>401,-8,401,-6</points>
<connection>
<GID>268</GID>
<name>SEL_1</name></connection>
<intersection>-6 13</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>380,33.5,380,36</points>
<connection>
<GID>368</GID>
<name>SEL_1</name></connection>
<intersection>36 20</intersection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>338.5,104,338.5,110.5</points>
<connection>
<GID>365</GID>
<name>SEL_1</name></connection>
<intersection>110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227.5,110.5,418.5,110.5</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>338.5 0</intersection>
<intersection>418.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>418.5,-39,418.5,110.5</points>
<connection>
<GID>262</GID>
<name>SEL_1</name></connection>
<intersection>-25 14</intersection>
<intersection>62.5 8</intersection>
<intersection>110.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>391,62.5,418.5,62.5</points>
<intersection>391 9</intersection>
<intersection>418.5 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>391,62.5,391,87</points>
<intersection>62.5 8</intersection>
<intersection>87 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>352,87,395.5,87</points>
<intersection>352 16</intersection>
<intersection>391 9</intersection>
<intersection>395.5 17</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>412,-25,418.5,-25</points>
<intersection>412 15</intersection>
<intersection>418.5 6</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>412,-28.5,412,-25</points>
<connection>
<GID>272</GID>
<name>SEL_1</name></connection>
<intersection>-25 14</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>352,86,352,87</points>
<connection>
<GID>241</GID>
<name>SEL_1</name></connection>
<intersection>87 10</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>395.5,2.5,395.5,87</points>
<connection>
<GID>266</GID>
<name>SEL_1</name></connection>
<intersection>25 24</intersection>
<intersection>46.5 22</intersection>
<intersection>68 19</intersection>
<intersection>87 10</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>364,68,395.5,68</points>
<intersection>364 20</intersection>
<intersection>395.5 17</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>364,65,364,68</points>
<connection>
<GID>360</GID>
<name>SEL_1</name></connection>
<intersection>68 19</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>374.5,46.5,395.5,46.5</points>
<intersection>374.5 25</intersection>
<intersection>395.5 17</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>385.5,25,395.5,25</points>
<intersection>385.5 26</intersection>
<intersection>395.5 17</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>374.5,43.5,374.5,46.5</points>
<connection>
<GID>366</GID>
<name>SEL_1</name></connection>
<intersection>46.5 22</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>385.5,23,385.5,25</points>
<connection>
<GID>369</GID>
<name>SEL_1</name></connection>
<intersection>25 24</intersection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203.5,-18,207,-18</points>
<connection>
<GID>371</GID>
<name>OUT_0</name></connection>
<intersection>207 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>207,-18,207,-12</points>
<intersection>-18 1</intersection>
<intersection>-12 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>207,-12,209,-12</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<intersection>207 7</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-24,208,-13</points>
<intersection>-24 3</intersection>
<intersection>-13 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>198,-24,208,-24</points>
<intersection>198 6</intersection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>208,-13,209,-13</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>208 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>198,-24,198,-23.5</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>-24 3</intersection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216.5,61,284,61</points>
<connection>
<GID>189</GID>
<name>load</name></connection>
<intersection>216.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>216.5,-10,216.5,61</points>
<intersection>-10 7</intersection>
<intersection>61 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>215,-10,216.5,-10</points>
<connection>
<GID>383</GID>
<name>OUT_3</name></connection>
<intersection>216.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,42.5,-34,42.5</points>
<connection>
<GID>118</GID>
<name>OUT_1</name></connection>
<connection>
<GID>148</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,41.5,-34,41.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-43.5,51,-43.5,53</points>
<intersection>51 5</intersection>
<intersection>53 11</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-46.5,51,-43.5,51</points>
<intersection>-46.5 7</intersection>
<intersection>-43.5 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-46.5,50.5,-46.5,51</points>
<connection>
<GID>118</GID>
<name>load</name></connection>
<intersection>51 5</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-44,53,-43.5,53</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-43.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,40,36.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_10</name></connection>
<intersection>40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,40,39,40</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-11,218.5,37</points>
<intersection>-11 1</intersection>
<intersection>37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215,-11,218.5,-11</points>
<connection>
<GID>383</GID>
<name>OUT_2</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>218.5,37,285.5,37</points>
<connection>
<GID>232</GID>
<name>load</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>13,134.5,14,134.5</points>
<connection>
<GID>128</GID>
<name>OUT_7</name></connection>
<connection>
<GID>129</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>13,133.5,14,133.5</points>
<connection>
<GID>128</GID>
<name>OUT_6</name></connection>
<connection>
<GID>129</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>13,132.5,14,132.5</points>
<connection>
<GID>128</GID>
<name>OUT_5</name></connection>
<connection>
<GID>129</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>13,131.5,14,131.5</points>
<connection>
<GID>128</GID>
<name>OUT_4</name></connection>
<connection>
<GID>129</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>13,130.5,14,130.5</points>
<connection>
<GID>128</GID>
<name>OUT_3</name></connection>
<connection>
<GID>129</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>13,129.5,14,129.5</points>
<connection>
<GID>128</GID>
<name>OUT_2</name></connection>
<connection>
<GID>129</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>13,128.5,14,128.5</points>
<connection>
<GID>128</GID>
<name>OUT_1</name></connection>
<connection>
<GID>129</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>13,127.5,14,127.5</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>10,121.5,10,125.5</points>
<connection>
<GID>128</GID>
<name>clear</name></connection>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>26</ID>
<points>5.5,136.5,5.5,144</points>
<intersection>136.5 46</intersection>
<intersection>144 44</intersection></vsegment>
<hsegment>
<ID>44</ID>
<points>1,144,5.5,144</points>
<intersection>1 45</intersection>
<intersection>5.5 26</intersection></hsegment>
<vsegment>
<ID>45</ID>
<points>1,144,1,146</points>
<intersection>144 44</intersection>
<intersection>146 48</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>5.5,136.5,8,136.5</points>
<connection>
<GID>128</GID>
<name>load</name></connection>
<intersection>5.5 26</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>1,146,1,146</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>1 45</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71,61,-71,67.5</points>
<intersection>61 1</intersection>
<intersection>67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71,61,-68,61</points>
<connection>
<GID>147</GID>
<name>ADDRESS_7</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,67.5,-71,67.5</points>
<intersection>-97 3</intersection>
<intersection>-71 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-97,67.5,-97,70.5</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>67.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72,60,-72,65</points>
<intersection>60 1</intersection>
<intersection>65 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72,60,-68,60</points>
<connection>
<GID>147</GID>
<name>ADDRESS_6</name></connection>
<intersection>-72 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-97,65,-72,65</points>
<intersection>-97 4</intersection>
<intersection>-72 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-97,65,-97,66.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>65 3</intersection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73,59,-73,63</points>
<intersection>59 1</intersection>
<intersection>63 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,59,-68,59</points>
<connection>
<GID>147</GID>
<name>ADDRESS_5</name></connection>
<intersection>-73 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-97,63,-73,63</points>
<intersection>-97 4</intersection>
<intersection>-73 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-97,63,-97,63.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>63 3</intersection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74,58,-74,61</points>
<intersection>58 1</intersection>
<intersection>61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74,58,-68,58</points>
<connection>
<GID>147</GID>
<name>ADDRESS_4</name></connection>
<intersection>-74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,61,-74,61</points>
<intersection>-97 3</intersection>
<intersection>-74 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-97,60.5,-97,61</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>61 2</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74,54,-74,57</points>
<intersection>54 3</intersection>
<intersection>57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74,57,-68,57</points>
<connection>
<GID>147</GID>
<name>ADDRESS_3</name></connection>
<intersection>-74 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-97,54,-74,54</points>
<intersection>-97 4</intersection>
<intersection>-74 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-97,54,-97,57</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>54 3</intersection></vsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73,52,-73,56</points>
<intersection>52 2</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,56,-68,56</points>
<connection>
<GID>147</GID>
<name>ADDRESS_2</name></connection>
<intersection>-73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,52,-73,52</points>
<intersection>-97 3</intersection>
<intersection>-73 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-97,52,-97,53.5</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>52 2</intersection></vsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72,50,-72,55</points>
<intersection>50 2</intersection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72,55,-68,55</points>
<connection>
<GID>147</GID>
<name>ADDRESS_1</name></connection>
<intersection>-72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,50,-72,50</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>-72 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71,48,-71,54</points>
<intersection>48 2</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71,54,-68,54</points>
<connection>
<GID>147</GID>
<name>ADDRESS_0</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,48,-71,48</points>
<intersection>-97 3</intersection>
<intersection>-71 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-97,46.5,-97,48</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></vsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,112,96,119</points>
<intersection>112 2</intersection>
<intersection>119 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>96,112,97,112</points>
<connection>
<GID>154</GID>
<name>IN_7</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>92,119,96,119</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,111,95,116</points>
<intersection>111 1</intersection>
<intersection>116 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,111,97,111</points>
<connection>
<GID>154</GID>
<name>IN_6</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,116,95,116</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,110,94,113</points>
<intersection>110 1</intersection>
<intersection>113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,110,97,110</points>
<connection>
<GID>154</GID>
<name>IN_5</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,113,94,113</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>93,109,93,110</points>
<intersection>109 8</intersection>
<intersection>110 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>93,109,97,109</points>
<connection>
<GID>154</GID>
<name>IN_4</name></connection>
<intersection>93 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>92,110,93,110</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>93 7</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,107,93,108</points>
<intersection>107 2</intersection>
<intersection>108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,108,97,108</points>
<connection>
<GID>154</GID>
<name>IN_3</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,107,93,107</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92,104,94,104</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>94 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>94,104,94,107</points>
<intersection>104 1</intersection>
<intersection>107 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>94,107,97,107</points>
<connection>
<GID>154</GID>
<name>IN_2</name></connection>
<intersection>94 3</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,101,95,106</points>
<intersection>101 2</intersection>
<intersection>106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,106,97,106</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,101,95,101</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,98,96,105</points>
<intersection>98 2</intersection>
<intersection>105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,105,97,105</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,98,96,98</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,115,96.5,124.5</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>115 2</intersection>
<intersection>116 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>100,114,100,115</points>
<connection>
<GID>154</GID>
<name>load</name></connection>
<intersection>115 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>96.5,115,100,115</points>
<intersection>96.5 0</intersection>
<intersection>100 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>96.5,116,98,116</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,109,106,133.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,109,127,109</points>
<connection>
<GID>154</GID>
<name>OUT_4</name></connection>
<connection>
<GID>167</GID>
<name>IN_4</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,110,107,133.5</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,110,127,110</points>
<connection>
<GID>154</GID>
<name>OUT_5</name></connection>
<connection>
<GID>167</GID>
<name>IN_5</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,111,108,133.5</points>
<connection>
<GID>177</GID>
<name>IN_2</name></connection>
<intersection>111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,111,127,111</points>
<connection>
<GID>154</GID>
<name>OUT_6</name></connection>
<connection>
<GID>167</GID>
<name>IN_6</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,112,109,133.5</points>
<connection>
<GID>177</GID>
<name>IN_3</name></connection>
<intersection>112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,112,127,112</points>
<connection>
<GID>154</GID>
<name>OUT_7</name></connection>
<connection>
<GID>167</GID>
<name>IN_7</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,108,126,133.5</points>
<connection>
<GID>178</GID>
<name>IN_3</name></connection>
<intersection>108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,108,127,108</points>
<connection>
<GID>154</GID>
<name>OUT_3</name></connection>
<connection>
<GID>167</GID>
<name>IN_3</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,105,123,133.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,105,127,105</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,106,127,106</points>
<connection>
<GID>154</GID>
<name>OUT_1</name></connection>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<intersection>124 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>124,106,124,133.5</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>106 1</intersection></vsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,107,125,133.5</points>
<connection>
<GID>178</GID>
<name>IN_2</name></connection>
<intersection>107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,107,127,107</points>
<connection>
<GID>154</GID>
<name>OUT_2</name></connection>
<connection>
<GID>167</GID>
<name>IN_2</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>112,136.5,113,136.5</points>
<connection>
<GID>177</GID>
<name>carry_out</name></connection>
<connection>
<GID>178</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>95,136.5,96,136.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<connection>
<GID>177</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220.5,-12,220.5,12</points>
<intersection>-12 1</intersection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215,-12,220.5,-12</points>
<connection>
<GID>383</GID>
<name>OUT_1</name></connection>
<intersection>220.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,12,285,12</points>
<connection>
<GID>242</GID>
<name>load</name></connection>
<intersection>220.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,142.5,99.5,144.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>142.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>99.5,142.5,102.5,142.5</points>
<intersection>99.5 0</intersection>
<intersection>102.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102.5,141.5,102.5,142.5</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>142.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,141.5,103.5,143.5</points>
<connection>
<GID>177</GID>
<name>OUT_1</name></connection>
<intersection>143.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>102.5,143.5,102.5,144.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>143.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>102.5,143.5,103.5,143.5</points>
<intersection>102.5 1</intersection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,141.5,104.5,143.5</points>
<connection>
<GID>177</GID>
<name>OUT_2</name></connection>
<intersection>143.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104.5,143.5,105.5,143.5</points>
<intersection>104.5 0</intersection>
<intersection>105.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>105.5,143.5,105.5,144.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>143.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>105.5,142.5,108.5,142.5</points>
<intersection>105.5 4</intersection>
<intersection>108.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>105.5,141.5,105.5,142.5</points>
<connection>
<GID>177</GID>
<name>OUT_3</name></connection>
<intersection>142.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>108.5,142.5,108.5,144.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>142.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,143.5,119.5,144.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>143.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>120.5,141.5,120.5,143.5</points>
<connection>
<GID>178</GID>
<name>OUT_1</name></connection>
<intersection>143.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>119.5,143.5,120.5,143.5</points>
<intersection>119.5 0</intersection>
<intersection>120.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,141.5,121.5,143.5</points>
<connection>
<GID>178</GID>
<name>OUT_2</name></connection>
<intersection>143.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>121.5,143.5,122.5,143.5</points>
<intersection>121.5 0</intersection>
<intersection>122.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>122.5,143.5,122.5,144.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>143.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>122.5,141.5,122.5,142.5</points>
<connection>
<GID>178</GID>
<name>OUT_3</name></connection>
<intersection>142.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>122.5,142.5,125.5,142.5</points>
<intersection>122.5 1</intersection>
<intersection>125.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>125.5,142.5,125.5,144.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>142.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>119.5,141.5,119.5,142.5</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>142.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>116.5,142.5,119.5,142.5</points>
<intersection>116.5 3</intersection>
<intersection>119.5 1</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,142.5,116.5,144.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>142.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,28,-59.5,50.5</points>
<connection>
<GID>147</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>147</GID>
<name>DATA_IN_0</name></connection>
<intersection>28 17</intersection>
<intersection>41.5 28</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-68,28,-59.5,28</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-59.5,41.5,-49.5,41.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,29,-60.5,50.5</points>
<connection>
<GID>147</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>147</GID>
<name>DATA_IN_1</name></connection>
<intersection>29 17</intersection>
<intersection>42.5 46</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-68,29,-60.5,29</points>
<connection>
<GID>183</GID>
<name>OUT_1</name></connection>
<intersection>-60.5 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>-60.5,42.5,-49.5,42.5</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>-60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,30,-61.5,50.5</points>
<connection>
<GID>147</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>147</GID>
<name>DATA_IN_2</name></connection>
<intersection>30 10</intersection>
<intersection>43.5 38</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-68,30,-61.5,30</points>
<connection>
<GID>183</GID>
<name>OUT_2</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>-61.5,43.5,-49.5,43.5</points>
<connection>
<GID>118</GID>
<name>IN_2</name></connection>
<intersection>-61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-62.5,31,-62.5,50.5</points>
<connection>
<GID>147</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>147</GID>
<name>DATA_IN_3</name></connection>
<intersection>31 20</intersection>
<intersection>44.5 48</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-68,31,-62.5,31</points>
<connection>
<GID>183</GID>
<name>OUT_3</name></connection>
<intersection>-62.5 3</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>-62.5,44.5,-49.5,44.5</points>
<connection>
<GID>118</GID>
<name>IN_3</name></connection>
<intersection>-62.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,32,-63.5,50.5</points>
<connection>
<GID>147</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>147</GID>
<name>DATA_IN_4</name></connection>
<intersection>32 17</intersection>
<intersection>45.5 45</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-68,32,-63.5,32</points>
<connection>
<GID>183</GID>
<name>OUT_4</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-63.5,45.5,-49.5,45.5</points>
<connection>
<GID>118</GID>
<name>IN_4</name></connection>
<intersection>-63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,33,-64.5,50.5</points>
<connection>
<GID>147</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>147</GID>
<name>DATA_IN_5</name></connection>
<intersection>33 17</intersection>
<intersection>46.5 31</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-68,33,-64.5,33</points>
<connection>
<GID>183</GID>
<name>OUT_5</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>-64.5,46.5,-49.5,46.5</points>
<connection>
<GID>118</GID>
<name>IN_5</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,34,-65.5,50.5</points>
<connection>
<GID>147</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>147</GID>
<name>DATA_IN_6</name></connection>
<intersection>34 46</intersection>
<intersection>47.5 31</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>-65.5,47.5,-49.5,47.5</points>
<connection>
<GID>118</GID>
<name>IN_6</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>46</ID>
<points>-68,34,-65.5,34</points>
<connection>
<GID>183</GID>
<name>OUT_6</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,35,-66.5,50.5</points>
<connection>
<GID>147</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>147</GID>
<name>DATA_IN_7</name></connection>
<intersection>35 10</intersection>
<intersection>48.5 24</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-68,35,-66.5,35</points>
<connection>
<GID>183</GID>
<name>OUT_7</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-66.5,48.5,-49.5,48.5</points>
<connection>
<GID>118</GID>
<name>IN_7</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,49.5,-57,68</points>
<intersection>49.5 3</intersection>
<intersection>58 2</intersection>
<intersection>68 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-58,58,-57,58</points>
<connection>
<GID>147</GID>
<name>write_enable</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-70,49.5,-57,49.5</points>
<intersection>-70 4</intersection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-70,36.5,-70,49.5</points>
<connection>
<GID>183</GID>
<name>ENABLE_0</name></connection>
<intersection>49.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-59,68,-57,68</points>
<intersection>-59 6</intersection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-59,68,-59,69.5</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>68 5</intersection></vsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97.5,41,-73,41</points>
<intersection>-97.5 9</intersection>
<intersection>-73 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-73,35,-73,41</points>
<intersection>35 6</intersection>
<intersection>41 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-73,35,-72,35</points>
<connection>
<GID>183</GID>
<name>IN_7</name></connection>
<intersection>-73 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-97.5,41,-97.5,42</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-13,285,-13</points>
<connection>
<GID>244</GID>
<name>load</name></connection>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339.5,104,339.5,106</points>
<connection>
<GID>365</GID>
<name>SEL_0</name></connection>
<intersection>106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227.5,106,419.5,106</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>339.5 0</intersection>
<intersection>419.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>419.5,-39,419.5,106</points>
<connection>
<GID>262</GID>
<name>SEL_0</name></connection>
<intersection>-26 13</intersection>
<intersection>59.5 7</intersection>
<intersection>106 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>395,59.5,419.5,59.5</points>
<intersection>395 8</intersection>
<intersection>419.5 5</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>395,59.5,395,86</points>
<intersection>59.5 7</intersection>
<intersection>86 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>353,86,396.5,86</points>
<connection>
<GID>241</GID>
<name>SEL_0</name></connection>
<intersection>395 8</intersection>
<intersection>396.5 15</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>413,-26,419.5,-26</points>
<intersection>413 14</intersection>
<intersection>419.5 5</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>413,-28.5,413,-26</points>
<connection>
<GID>272</GID>
<name>SEL_0</name></connection>
<intersection>-26 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>396.5,2.5,396.5,86</points>
<connection>
<GID>266</GID>
<name>SEL_0</name></connection>
<intersection>24 20</intersection>
<intersection>45 16</intersection>
<intersection>66.5 17</intersection>
<intersection>86 9</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>375.5,45,396.5,45</points>
<intersection>375.5 21</intersection>
<intersection>396.5 15</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>365,66.5,396.5,66.5</points>
<intersection>365 18</intersection>
<intersection>396.5 15</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>365,65,365,66.5</points>
<connection>
<GID>360</GID>
<name>SEL_0</name></connection>
<intersection>66.5 17</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>386.5,24,396.5,24</points>
<intersection>386.5 22</intersection>
<intersection>396.5 15</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>375.5,43.5,375.5,45</points>
<connection>
<GID>366</GID>
<name>SEL_0</name></connection>
<intersection>45 16</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>386.5,23,386.5,24</points>
<connection>
<GID>369</GID>
<name>SEL_0</name></connection>
<intersection>24 20</intersection></vsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>406.5,58,479,58</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>406.5 8</intersection>
<intersection>460.5 11</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>406.5,58,406.5,99</points>
<intersection>58 1</intersection>
<intersection>99 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>341.5,99,406.5,99</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<intersection>406.5 8</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>460.5,55.5,460.5,58</points>
<connection>
<GID>258</GID>
<name>IN_7</name></connection>
<intersection>58 1</intersection></vsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200.5,58,281,58</points>
<connection>
<GID>189</GID>
<name>IN_6</name></connection>
<intersection>200.5 15</intersection>
<intersection>234.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>234.5,34,234.5,58</points>
<intersection>34 6</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>234.5,34,282.5,34</points>
<connection>
<GID>232</GID>
<name>IN_6</name></connection>
<intersection>234.5 5</intersection>
<intersection>250.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>250.5,9,250.5,34</points>
<intersection>9 9</intersection>
<intersection>34 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>250.5,9,282,9</points>
<connection>
<GID>242</GID>
<name>IN_6</name></connection>
<intersection>250.5 8</intersection>
<intersection>266.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>266.5,-16,266.5,9</points>
<intersection>-16 11</intersection>
<intersection>9 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>266.5,-16,282,-16</points>
<connection>
<GID>244</GID>
<name>IN_6</name></connection>
<intersection>266.5 10</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>200.5,52.5,200.5,58</points>
<intersection>52.5 16</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>191,52.5,200.5,52.5</points>
<intersection>191 20</intersection>
<intersection>200.5 15</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>191,41.5,191,52.5</points>
<intersection>41.5 22</intersection>
<intersection>52.5 16</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>189.5,41.5,191,41.5</points>
<connection>
<GID>95</GID>
<name>OUT_6</name></connection>
<intersection>191 20</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-74,24,-74,29</points>
<intersection>24 6</intersection>
<intersection>29 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-74,29,-72,29</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>-74 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-97.5,24,-74,24</points>
<intersection>-97.5 9</intersection>
<intersection>-74 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-97.5,21.5,-97.5,24</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>24 6</intersection></vsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,18,-84.5,28</points>
<intersection>18 11</intersection>
<intersection>28 12</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-97.5,18,-84.5,18</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-84.5,28,-72,28</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<hsegment>
<ID>18</ID>
<points>-30,48.5,-14.5,48.5</points>
<connection>
<GID>148</GID>
<name>OUT_7</name></connection>
<connection>
<GID>273</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>-16.5,46,-16.5,47.5</points>
<intersection>46 18</intersection>
<intersection>47.5 19</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-16.5,46,-15.5,46</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>-16.5 11</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-30,47.5,-16.5,47.5</points>
<connection>
<GID>148</GID>
<name>OUT_6</name></connection>
<intersection>-16.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>-17,43.5,-17,46.5</points>
<intersection>43.5 12</intersection>
<intersection>46.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-17,43.5,-15.5,43.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>-17 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-30,46.5,-17,46.5</points>
<connection>
<GID>148</GID>
<name>OUT_5</name></connection>
<intersection>-17 11</intersection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>-18,41,-18,45.5</points>
<intersection>41 12</intersection>
<intersection>45.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-18,41,-15.5,41</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-18 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-30,45.5,-18,45.5</points>
<connection>
<GID>148</GID>
<name>OUT_4</name></connection>
<intersection>-18 11</intersection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>-18.5,38,-18.5,44.5</points>
<intersection>38 13</intersection>
<intersection>44.5 14</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-18.5,38,-15.5,38</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>-18.5 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-30,44.5,-18.5,44.5</points>
<connection>
<GID>148</GID>
<name>OUT_3</name></connection>
<intersection>-18.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>-19,35,-19,43.5</points>
<intersection>35 12</intersection>
<intersection>43.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-19,35,-15,35</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>-19 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-30,43.5,-19,43.5</points>
<connection>
<GID>148</GID>
<name>OUT_2</name></connection>
<intersection>-19 11</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>-19.5,32,-19.5,42.5</points>
<intersection>32 12</intersection>
<intersection>42.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-19.5,32,-15,32</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>-19.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-30,42.5,-19.5,42.5</points>
<connection>
<GID>148</GID>
<name>OUT_1</name></connection>
<intersection>-19.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>14</ID>
<points>-20,29,-20,41.5</points>
<intersection>29 15</intersection>
<intersection>41.5 16</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-20,29,-15,29</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>-20 14</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-30,41.5,-20,41.5</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>-20 14</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,135.5,-62.5,137.5</points>
<connection>
<GID>214</GID>
<name>load</name></connection>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-60.5,123,-60.5,124.5</points>
<connection>
<GID>214</GID>
<name>clear</name></connection>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73,114.5,-73,126.5</points>
<intersection>114.5 2</intersection>
<intersection>126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,126.5,-65.5,126.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,114.5,-73,114.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>-73 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74.5,118,-74.5,127.5</points>
<intersection>118 2</intersection>
<intersection>127.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74.5,127.5,-65.5,127.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>-74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,118,-74.5,118</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>-74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76,123,-76,128.5</points>
<intersection>123 2</intersection>
<intersection>128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,128.5,-65.5,128.5</points>
<connection>
<GID>214</GID>
<name>IN_2</name></connection>
<intersection>-76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,123,-76,123</points>
<intersection>-79.5 3</intersection>
<intersection>-76 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-79.5,121.5,-79.5,123</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>123 2</intersection></vsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,125,-78,129.5</points>
<intersection>125 2</intersection>
<intersection>129.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-78,129.5,-65.5,129.5</points>
<connection>
<GID>214</GID>
<name>IN_3</name></connection>
<intersection>-78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,125,-78,125</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>-78 0</intersection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,130.5,-65.5,130.5</points>
<connection>
<GID>214</GID>
<name>IN_4</name></connection>
<intersection>-79.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-79.5,128.5,-79.5,130.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>130.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,131.5,-65.5,131.5</points>
<connection>
<GID>214</GID>
<name>IN_5</name></connection>
<connection>
<GID>226</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75.5,132.5,-75.5,135</points>
<intersection>132.5 1</intersection>
<intersection>135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75.5,132.5,-65.5,132.5</points>
<connection>
<GID>214</GID>
<name>IN_6</name></connection>
<intersection>-75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,135,-75.5,135</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>-75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72,133.5,-72,138.5</points>
<intersection>133.5 3</intersection>
<intersection>138.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,138.5,-72,138.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>-72 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-72,133.5,-65.5,133.5</points>
<connection>
<GID>214</GID>
<name>IN_7</name></connection>
<intersection>-72 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,133.5,-57.5,140</points>
<connection>
<GID>214</GID>
<name>OUT_7</name></connection>
<intersection>140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57.5,140,-49,140</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,132.5,-54,137.5</points>
<intersection>132.5 2</intersection>
<intersection>137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,137.5,-49,137.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>-54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,132.5,-54,132.5</points>
<connection>
<GID>214</GID>
<name>OUT_6</name></connection>
<intersection>-54 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,131.5,-52,135</points>
<intersection>131.5 2</intersection>
<intersection>135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52,135,-49,135</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>-52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,131.5,-52,131.5</points>
<connection>
<GID>214</GID>
<name>OUT_5</name></connection>
<intersection>-52 0</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51,130.5,-51,132</points>
<intersection>130.5 2</intersection>
<intersection>132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51,132,-49,132</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>-51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,130.5,-51,130.5</points>
<connection>
<GID>214</GID>
<name>OUT_4</name></connection>
<intersection>-51 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-57.5,129.5,-49,129.5</points>
<connection>
<GID>214</GID>
<name>OUT_3</name></connection>
<connection>
<GID>237</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,126,-54.5,128.5</points>
<intersection>126 1</intersection>
<intersection>128.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54.5,126,-49,126</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,128.5,-54.5,128.5</points>
<connection>
<GID>214</GID>
<name>OUT_2</name></connection>
<intersection>-54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,123,-55.5,127.5</points>
<intersection>123 1</intersection>
<intersection>127.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55.5,123,-49,123</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>-55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,127.5,-55.5,127.5</points>
<connection>
<GID>214</GID>
<name>OUT_1</name></connection>
<intersection>-55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,120,-56.5,126.5</points>
<intersection>120 1</intersection>
<intersection>126.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56.5,120,-49,120</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,126.5,-56.5,126.5</points>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203,57,281,57</points>
<connection>
<GID>189</GID>
<name>IN_5</name></connection>
<intersection>203 10</intersection>
<intersection>232.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>232.5,33,232.5,57</points>
<intersection>33 9</intersection>
<intersection>57 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>232.5,33,282.5,33</points>
<connection>
<GID>232</GID>
<name>IN_5</name></connection>
<intersection>232.5 8</intersection>
<intersection>248.5 12</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>203,47.5,203,57</points>
<intersection>47.5 11</intersection>
<intersection>57 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>192,47.5,203,47.5</points>
<intersection>192 19</intersection>
<intersection>203 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>248.5,8,248.5,33</points>
<intersection>8 13</intersection>
<intersection>33 9</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>248.5,8,282,8</points>
<connection>
<GID>242</GID>
<name>IN_5</name></connection>
<intersection>248.5 12</intersection>
<intersection>264.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>264.5,-17,264.5,8</points>
<intersection>-17 15</intersection>
<intersection>8 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>264.5,-17,282,-17</points>
<connection>
<GID>244</GID>
<name>IN_5</name></connection>
<intersection>264.5 14</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>192,40.5,192,47.5</points>
<intersection>40.5 21</intersection>
<intersection>47.5 11</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>189.5,40.5,192,40.5</points>
<connection>
<GID>95</GID>
<name>OUT_5</name></connection>
<intersection>192 19</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,56,281,56</points>
<connection>
<GID>189</GID>
<name>IN_4</name></connection>
<intersection>205 7</intersection>
<intersection>230.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>230.5,32,230.5,56</points>
<intersection>32 6</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>230.5,32,282.5,32</points>
<connection>
<GID>232</GID>
<name>IN_4</name></connection>
<intersection>230.5 5</intersection>
<intersection>246.5 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>205,45,205,56</points>
<intersection>45 8</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>193,45,205,45</points>
<intersection>193 16</intersection>
<intersection>205 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>246.5,7,246.5,32</points>
<intersection>7 10</intersection>
<intersection>32 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>246.5,7,282,7</points>
<connection>
<GID>242</GID>
<name>IN_4</name></connection>
<intersection>246.5 9</intersection>
<intersection>262.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>262.5,-18,262.5,7</points>
<intersection>-18 12</intersection>
<intersection>7 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>262.5,-18,282,-18</points>
<connection>
<GID>244</GID>
<name>IN_4</name></connection>
<intersection>262.5 11</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>193,39.5,193,45</points>
<intersection>39.5 17</intersection>
<intersection>45 8</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>189.5,39.5,193,39.5</points>
<connection>
<GID>95</GID>
<name>OUT_4</name></connection>
<intersection>193 16</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207.5,55,281,55</points>
<connection>
<GID>189</GID>
<name>IN_3</name></connection>
<intersection>207.5 7</intersection>
<intersection>228.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>228.5,31,228.5,55</points>
<intersection>31 6</intersection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>228.5,31,282.5,31</points>
<connection>
<GID>232</GID>
<name>IN_3</name></connection>
<intersection>228.5 5</intersection>
<intersection>244.5 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>207.5,41.5,207.5,55</points>
<intersection>41.5 8</intersection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>194,41.5,207.5,41.5</points>
<intersection>194 14</intersection>
<intersection>207.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>244.5,6,244.5,31</points>
<intersection>6 10</intersection>
<intersection>31 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>244.5,6,282,6</points>
<connection>
<GID>242</GID>
<name>IN_3</name></connection>
<intersection>244.5 9</intersection>
<intersection>260.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>260.5,-19,260.5,6</points>
<intersection>-19 12</intersection>
<intersection>6 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>260.5,-19,282,-19</points>
<connection>
<GID>244</GID>
<name>IN_3</name></connection>
<intersection>260.5 11</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>194,38.5,194,41.5</points>
<intersection>38.5 15</intersection>
<intersection>41.5 8</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>189.5,38.5,194,38.5</points>
<connection>
<GID>95</GID>
<name>OUT_3</name></connection>
<intersection>194 14</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209.5,54,281,54</points>
<connection>
<GID>189</GID>
<name>IN_2</name></connection>
<intersection>209.5 7</intersection>
<intersection>226.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>226.5,30,226.5,54</points>
<intersection>30 6</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>226.5,30,282.5,30</points>
<connection>
<GID>232</GID>
<name>IN_2</name></connection>
<intersection>226.5 5</intersection>
<intersection>242.5 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>209.5,40.5,209.5,54</points>
<intersection>40.5 8</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>197,40.5,209.5,40.5</points>
<intersection>197 14</intersection>
<intersection>209.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>242.5,5,242.5,30</points>
<intersection>5 10</intersection>
<intersection>30 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>242.5,5,282,5</points>
<connection>
<GID>242</GID>
<name>IN_2</name></connection>
<intersection>242.5 9</intersection>
<intersection>258.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>258.5,-20,258.5,5</points>
<intersection>-20 12</intersection>
<intersection>5 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>258.5,-20,282,-20</points>
<connection>
<GID>244</GID>
<name>IN_2</name></connection>
<intersection>258.5 11</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>197,37.5,197,40.5</points>
<intersection>37.5 17</intersection>
<intersection>40.5 8</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>189.5,37.5,197,37.5</points>
<connection>
<GID>95</GID>
<name>OUT_2</name></connection>
<intersection>197 14</intersection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>211.5,53,281,53</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>211.5 7</intersection>
<intersection>224.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>224.5,29,224.5,53</points>
<intersection>29 6</intersection>
<intersection>53 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>224.5,29,282.5,29</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<intersection>224.5 5</intersection>
<intersection>240.5 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>211.5,36.5,211.5,53</points>
<intersection>36.5 8</intersection>
<intersection>53 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>189.5,36.5,211.5,36.5</points>
<connection>
<GID>95</GID>
<name>OUT_1</name></connection>
<intersection>211.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>240.5,4,240.5,29</points>
<intersection>4 10</intersection>
<intersection>29 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>240.5,4,282,4</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>240.5 9</intersection>
<intersection>256.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>256.5,-21,256.5,4</points>
<intersection>-21 12</intersection>
<intersection>4 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>256.5,-21,282,-21</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>256.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222.5,52,281,52</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>222.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>222.5,28,222.5,52</points>
<intersection>28 6</intersection>
<intersection>30 16</intersection>
<intersection>52 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>222.5,28,282.5,28</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>222.5 5</intersection>
<intersection>238.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>238.5,3,238.5,28</points>
<intersection>3 10</intersection>
<intersection>28 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>238.5,3,282,3</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>238.5 9</intersection>
<intersection>254.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>254.5,-22,254.5,3</points>
<intersection>-22 12</intersection>
<intersection>3 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>254.5,-22,282,-22</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>254.5 11</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>201.5,30,222.5,30</points>
<intersection>201.5 17</intersection>
<intersection>222.5 5</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>201.5,30,201.5,35.5</points>
<intersection>30 16</intersection>
<intersection>35.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>189.5,35.5,201.5,35.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>201.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,134.5,3,141.5</points>
<intersection>134.5 2</intersection>
<intersection>141.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,141.5,3,141.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,134.5,5,134.5</points>
<connection>
<GID>128</GID>
<name>IN_7</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,133.5,1,138</points>
<intersection>133.5 1</intersection>
<intersection>138 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,133.5,5,133.5</points>
<connection>
<GID>128</GID>
<name>IN_6</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,138,1,138</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,132.5,5,132.5</points>
<connection>
<GID>128</GID>
<name>IN_5</name></connection>
<intersection>-0.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-0.5,132.5,-0.5,134.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>132.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,131.5,5,131.5</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,128,1,130.5</points>
<intersection>128 2</intersection>
<intersection>130.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,130.5,5,130.5</points>
<connection>
<GID>128</GID>
<name>IN_3</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,128,1,128</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,124.5,2,129.5</points>
<intersection>124.5 2</intersection>
<intersection>129.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,129.5,5,129.5</points>
<connection>
<GID>128</GID>
<name>IN_2</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,124.5,2,124.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,121,3,128.5</points>
<intersection>121 2</intersection>
<intersection>128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,128.5,5,128.5</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,121,3,121</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,117.5,2,127.5</points>
<intersection>117.5 7</intersection>
<intersection>127.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-0.5,117.5,2,117.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>2,127.5,5,127.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189.5,59,281,59</points>
<connection>
<GID>189</GID>
<name>IN_7</name></connection>
<intersection>189.5 20</intersection>
<intersection>236.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>236.5,35,236.5,59</points>
<intersection>35 4</intersection>
<intersection>59 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>236.5,35,282.5,35</points>
<connection>
<GID>232</GID>
<name>IN_7</name></connection>
<intersection>236.5 3</intersection>
<intersection>252.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>252.5,10,252.5,35</points>
<intersection>10 6</intersection>
<intersection>35 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>252.5,10,282,10</points>
<connection>
<GID>242</GID>
<name>IN_7</name></connection>
<intersection>252.5 5</intersection>
<intersection>268.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>268.5,-15,268.5,10</points>
<intersection>-15 8</intersection>
<intersection>10 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>268.5,-15,282,-15</points>
<connection>
<GID>244</GID>
<name>IN_7</name></connection>
<intersection>268.5 7</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>189.5,42.5,189.5,59</points>
<connection>
<GID>95</GID>
<name>OUT_7</name></connection>
<intersection>59 1</intersection></vsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,20,408.5,89.5</points>
<intersection>20 1</intersection>
<intersection>89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,20,481,20</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection>
<intersection>462.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>347.5,89.5,408.5,89.5</points>
<connection>
<GID>385</GID>
<name>OUT</name></connection>
<intersection>408.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>462.5,17.5,462.5,20</points>
<connection>
<GID>101</GID>
<name>IN_7</name></connection>
<intersection>20 1</intersection></vsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,95,-67,124.5</points>
<intersection>95 3</intersection>
<intersection>124.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-67,124.5,-62.5,124.5</points>
<connection>
<GID>214</GID>
<name>clock</name></connection>
<intersection>-67 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-67,95,100,95</points>
<intersection>-67 0</intersection>
<intersection>-21.5 6</intersection>
<intersection>-12.5 4</intersection>
<intersection>8 8</intersection>
<intersection>100 7</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12.5,59,-12.5,95</points>
<intersection>59 5</intersection>
<intersection>95 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-58,59,-12.5,59</points>
<connection>
<GID>147</GID>
<name>write_clock</name></connection>
<intersection>-37 9</intersection>
<intersection>-12.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-21.5,95,-21.5,100</points>
<connection>
<GID>343</GID>
<name>CLK</name></connection>
<intersection>95 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>100,-2,100,103</points>
<connection>
<GID>154</GID>
<name>clock</name></connection>
<intersection>-2 15</intersection>
<intersection>23 14</intersection>
<intersection>48 17</intersection>
<intersection>71.5 19</intersection>
<intersection>95 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>8,95,8,125.5</points>
<connection>
<GID>128</GID>
<name>clock</name></connection>
<intersection>95 3</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-37,39.5,-37,59</points>
<intersection>39.5 10</intersection>
<intersection>59 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-46.5,39.5,-37,39.5</points>
<connection>
<GID>118</GID>
<name>clock</name></connection>
<intersection>-37 9</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>100,23,285,23</points>
<intersection>100 7</intersection>
<intersection>285 24</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>100,-2,285,-2</points>
<intersection>100 7</intersection>
<intersection>285 24</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>100,48,285.5,48</points>
<intersection>100 7</intersection>
<intersection>285.5 23</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>100,71.5,284,71.5</points>
<intersection>100 7</intersection>
<intersection>284 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>284,50,284,71.5</points>
<connection>
<GID>189</GID>
<name>clock</name></connection>
<intersection>71.5 19</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>285.5,26,285.5,48</points>
<connection>
<GID>232</GID>
<name>clock</name></connection>
<intersection>48 17</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>285,-24,285,23</points>
<connection>
<GID>242</GID>
<name>clock</name></connection>
<connection>
<GID>244</GID>
<name>clock</name></connection>
<intersection>-2 15</intersection>
<intersection>23 14</intersection></vsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-85,34,-85,38</points>
<intersection>34 1</intersection>
<intersection>38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-85,34,-72,34</points>
<connection>
<GID>183</GID>
<name>IN_6</name></connection>
<intersection>-85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-98,38,-85,38</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>-85 0</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,33,-84.5,35</points>
<intersection>33 1</intersection>
<intersection>35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84.5,33,-72,33</points>
<connection>
<GID>183</GID>
<name>IN_5</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97.5,35,-84.5,35</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97.5,32,-72,32</points>
<connection>
<GID>183</GID>
<name>IN_4</name></connection>
<connection>
<GID>346</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290.5,84,349,84</points>
<connection>
<GID>241</GID>
<name>IN_3</name></connection>
<intersection>290.5 8</intersection>
<intersection>310.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>310.5,73,310.5,84</points>
<intersection>73 4</intersection>
<intersection>84 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>310.5,73,355,73</points>
<connection>
<GID>243</GID>
<name>IN_3</name></connection>
<intersection>310.5 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>290.5,58,290.5,84</points>
<intersection>58 9</intersection>
<intersection>84 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>289,58,290.5,58</points>
<connection>
<GID>189</GID>
<name>OUT_6</name></connection>
<intersection>290.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-91.5,30,-72,30</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>-91.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-91.5,25,-91.5,30</points>
<intersection>25 6</intersection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-97.5,25,-91.5,25</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>-91.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97.5,28.5,-72,28.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>-72 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-72,28.5,-72,31</points>
<connection>
<GID>183</GID>
<name>IN_3</name></connection>
<intersection>28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,98,133,105</points>
<intersection>98 1</intersection>
<intersection>105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,98,145.5,98</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,105,133,105</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,103,134,106</points>
<intersection>103 1</intersection>
<intersection>106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,103,145.5,103</points>
<intersection>134 0</intersection>
<intersection>145.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,106,134,106</points>
<connection>
<GID>167</GID>
<name>OUT_1</name></connection>
<intersection>134 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>145.5,101,145.5,103</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>103 1</intersection></vsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,113.5,132.5,124.5</points>
<intersection>113.5 2</intersection>
<intersection>124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,124.5,139,124.5</points>
<intersection>132.5 0</intersection>
<intersection>139 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129,113.5,132.5,113.5</points>
<connection>
<GID>167</GID>
<name>ENABLE_0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>139,124.5,139,128.5</points>
<intersection>124.5 1</intersection>
<intersection>128.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>139,128.5,139,128.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>139 5</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,104,135.5,107</points>
<intersection>104 2</intersection>
<intersection>107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,107,135.5,107</points>
<connection>
<GID>167</GID>
<name>OUT_2</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135.5,104,145.5,104</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,107,138,108</points>
<intersection>107 1</intersection>
<intersection>108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,107,145,107</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,108,138,108</points>
<connection>
<GID>167</GID>
<name>OUT_3</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,109,140,110</points>
<intersection>109 1</intersection>
<intersection>110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,109,140,109</points>
<connection>
<GID>167</GID>
<name>OUT_4</name></connection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140,110,145,110</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,110,139.5,112.5</points>
<intersection>110 2</intersection>
<intersection>112.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139.5,112.5,145,112.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,110,139.5,110</points>
<connection>
<GID>167</GID>
<name>OUT_5</name></connection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,111,138,115</points>
<intersection>111 1</intersection>
<intersection>115 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,111,138,111</points>
<connection>
<GID>167</GID>
<name>OUT_6</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,115,145,115</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,112,136.5,117.5</points>
<intersection>112 2</intersection>
<intersection>117.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,117.5,146,117.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,112,136.5,112</points>
<connection>
<GID>167</GID>
<name>OUT_7</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>297.5,82,349,82</points>
<connection>
<GID>241</GID>
<name>IN_2</name></connection>
<intersection>297.5 5</intersection>
<intersection>308.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>308.5,71,308.5,82</points>
<intersection>71 4</intersection>
<intersection>82 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>308.5,71,355,71</points>
<connection>
<GID>243</GID>
<name>IN_2</name></connection>
<intersection>308.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>297.5,34,297.5,82</points>
<intersection>34 6</intersection>
<intersection>82 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>290.5,34,297.5,34</points>
<connection>
<GID>232</GID>
<name>OUT_6</name></connection>
<intersection>297.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>299.5,9,299.5,80</points>
<intersection>9 1</intersection>
<intersection>80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,9,299.5,9</points>
<connection>
<GID>242</GID>
<name>OUT_6</name></connection>
<intersection>299.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>299.5,80,349,80</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<intersection>299.5 0</intersection>
<intersection>306.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>306.5,69,306.5,80</points>
<intersection>69 4</intersection>
<intersection>80 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>306.5,69,355,69</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>306.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,64.5,24,132.5</points>
<intersection>64.5 1</intersection>
<intersection>132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,64.5,30,64.5</points>
<connection>
<GID>364</GID>
<name>ADDRESS_3</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,132.5,24,132.5</points>
<connection>
<GID>129</GID>
<name>OUT_5</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-15,295.5,96</points>
<intersection>-15 1</intersection>
<intersection>96 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-15,295.5,-15</points>
<connection>
<GID>244</GID>
<name>OUT_7</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295.5,96,335.5,96</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection>
<intersection>297.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>297.5,86.5,297.5,96</points>
<intersection>86.5 4</intersection>
<intersection>96 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>297.5,86.5,341.5,86.5</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>297.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,21.5,31.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_15</name></connection>
<intersection>21.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31.5,21.5,32,21.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,25,32.5,56</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<connection>
<GID>364</GID>
<name>DATA_OUT_14</name></connection></vsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,33.5,34.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_12</name></connection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,33.5,34.5,33.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,29,33.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_13</name></connection>
<intersection>29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,29,34,29</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-16,302,78</points>
<intersection>-16 1</intersection>
<intersection>78 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-16,302,-16</points>
<connection>
<GID>244</GID>
<name>OUT_6</name></connection>
<intersection>302 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>302,78,349,78</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>302 0</intersection>
<intersection>304.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>304.5,67,304.5,78</points>
<intersection>67 4</intersection>
<intersection>78 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>304.5,67,355,67</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>304.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355,81,447.5,81</points>
<connection>
<GID>241</GID>
<name>OUT</name></connection>
<intersection>447.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>447.5,54.5,447.5,81</points>
<intersection>54.5 5</intersection>
<intersection>81 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>447.5,54.5,460.5,54.5</points>
<connection>
<GID>258</GID>
<name>IN_6</name></connection>
<intersection>447.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>407,22,407,70</points>
<intersection>22 1</intersection>
<intersection>70 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>407,22,478,22</points>
<intersection>407 0</intersection>
<intersection>461 4</intersection>
<intersection>478 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>361,70,407,70</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<intersection>407 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>478,17,478,22</points>
<intersection>17 6</intersection>
<intersection>22 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>461,16.5,461,22</points>
<intersection>16.5 5</intersection>
<intersection>22 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>461,16.5,462.5,16.5</points>
<connection>
<GID>101</GID>
<name>IN_6</name></connection>
<intersection>461 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>478,17,481,17</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>478 3</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-56.5,422.5,-56.5</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>290 6</intersection>
<intersection>414 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>414,-56.5,414,-47</points>
<intersection>-56.5 1</intersection>
<intersection>-47 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>414,-47,415.5,-47</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>414 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>290,-56.5,290,-22</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>335.5,-54.5,335.5,3</points>
<intersection>-54.5 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>335.5,-54.5,422.5,-54.5</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>335.5 0</intersection>
<intersection>412 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>290,3,335.5,3</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>335.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>412,-54.5,412,-45</points>
<intersection>-54.5 1</intersection>
<intersection>-45 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>412,-45,415.5,-45</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>412 3</intersection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,65.5,25,133.5</points>
<intersection>65.5 1</intersection>
<intersection>133.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,65.5,30,65.5</points>
<connection>
<GID>364</GID>
<name>ADDRESS_4</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,133.5,25,133.5</points>
<connection>
<GID>129</GID>
<name>OUT_6</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,66.5,26,134.5</points>
<intersection>66.5 1</intersection>
<intersection>134.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,66.5,30,66.5</points>
<connection>
<GID>364</GID>
<name>ADDRESS_5</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,134.5,26,134.5</points>
<connection>
<GID>129</GID>
<name>OUT_7</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,136,23,141.5</points>
<intersection>136 2</intersection>
<intersection>141.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>16,136,23,136</points>
<connection>
<GID>129</GID>
<name>ENABLE_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23,141.5,23,141.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,42.5,37.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_9</name></connection>
<intersection>42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,42.5,39,42.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,107.5,28.5,123</points>
<intersection>107.5 1</intersection>
<intersection>123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,107.5,37,107.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,123,28.5,123</points>
<intersection>18 3</intersection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,123,18,127.5</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></vsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,110.5,31,124</points>
<intersection>110.5 1</intersection>
<intersection>124 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,110.5,37,110.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,124,31,124</points>
<intersection>19 3</intersection>
<intersection>31 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,124,19,128.5</points>
<intersection>124 2</intersection>
<intersection>128.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>18,128.5,19,128.5</points>
<connection>
<GID>129</GID>
<name>OUT_1</name></connection>
<intersection>19 3</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,113.5,32,125.5</points>
<intersection>113.5 2</intersection>
<intersection>125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,125.5,32,125.5</points>
<intersection>20.5 3</intersection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,113.5,37,113.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,125.5,20.5,129.5</points>
<intersection>125.5 1</intersection>
<intersection>129.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>18,129.5,20.5,129.5</points>
<connection>
<GID>129</GID>
<name>OUT_2</name></connection>
<intersection>20.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,130.5,23,130.5</points>
<connection>
<GID>129</GID>
<name>OUT_3</name></connection>
<intersection>23 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,126.5,23,130.5</points>
<intersection>126.5 4</intersection>
<intersection>130.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>23,126.5,33.5,126.5</points>
<intersection>23 3</intersection>
<intersection>33.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>33.5,116.5,33.5,126.5</points>
<intersection>116.5 6</intersection>
<intersection>126.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>33.5,116.5,36.5,116.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>33.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,119.5,35,129</points>
<intersection>119.5 2</intersection>
<intersection>122 3</intersection>
<intersection>124.5 4</intersection>
<intersection>127 5</intersection>
<intersection>129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,129,35,129</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,119.5,36.5,119.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,122,36.5,122</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35,124.5,36.5,124.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>35,127,37.5,127</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,50,46.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_0</name></connection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,50,46.5,50</points>
<intersection>28.5 2</intersection>
<intersection>46.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>28.5,50,28.5,61.5</points>
<intersection>50 1</intersection>
<intersection>61.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>28.5,61.5,30,61.5</points>
<connection>
<GID>364</GID>
<name>ADDRESS_0</name></connection>
<intersection>28.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,50.5,45.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_1</name></connection>
<intersection>50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,50.5,45.5,50.5</points>
<intersection>27 2</intersection>
<intersection>45.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>27,50.5,27,62.5</points>
<intersection>50.5 1</intersection>
<intersection>62.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>27,62.5,30,62.5</points>
<connection>
<GID>364</GID>
<name>ADDRESS_1</name></connection>
<intersection>27 2</intersection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,52.5,25.5,63.5</points>
<intersection>52.5 2</intersection>
<intersection>63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,63.5,30,63.5</points>
<connection>
<GID>364</GID>
<name>ADDRESS_2</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,52.5,44.5,52.5</points>
<intersection>25.5 0</intersection>
<intersection>44.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44.5,52.5,44.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_2</name></connection>
<intersection>52.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,-10,180,66</points>
<intersection>-10 2</intersection>
<intersection>44 3</intersection>
<intersection>66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180,66,182,66</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>180,-10,209,-10</points>
<connection>
<GID>383</GID>
<name>ENABLE</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>180,44,187.5,44</points>
<connection>
<GID>95</GID>
<name>ENABLE_0</name></connection>
<intersection>180 0</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,45.5,38.5,56</points>
<connection>
<GID>364</GID>
<name>DATA_OUT_8</name></connection>
<intersection>45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,45.5,41.5,45.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>120,-67,120,-67</points>
<connection>
<GID>320</GID>
<name>carry_out</name></connection>
<connection>
<GID>321</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-80,100.5,-52</points>
<intersection>-80 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-80,117,-80</points>
<connection>
<GID>321</GID>
<name>IN_3</name></connection>
<intersection>100.5 0</intersection>
<intersection>117 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-52,100.5,-52</points>
<connection>
<GID>322</GID>
<name>OUT_3</name></connection>
<intersection>100.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117,-84.5,117,-80</points>
<intersection>-84.5 4</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>117,-84.5,117.5,-84.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>117 3</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-79,99.5,-54</points>
<intersection>-79 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-79,117,-79</points>
<connection>
<GID>321</GID>
<name>IN_2</name></connection>
<intersection>99.5 0</intersection>
<intersection>117 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-54,99.5,-54</points>
<connection>
<GID>322</GID>
<name>OUT_2</name></connection>
<intersection>99.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117,-90,117,-79</points>
<intersection>-90 4</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>117,-90,117.5,-90</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>117 3</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-78,98.5,-56</points>
<intersection>-78 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-78,117,-78</points>
<connection>
<GID>321</GID>
<name>IN_1</name></connection>
<intersection>98.5 0</intersection>
<intersection>116.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-56,98.5,-56</points>
<connection>
<GID>322</GID>
<name>OUT_1</name></connection>
<intersection>98.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,-95.5,116.5,-78</points>
<intersection>-95.5 4</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>116.5,-95.5,117.5,-95.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>116.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-77,97.5,-58</points>
<intersection>-77 1</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-77,117,-77</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>97.5 0</intersection>
<intersection>116.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-58,97.5,-58</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,-101,116.5,-77</points>
<intersection>-101 4</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>116.5,-101,117.5,-101</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>116.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-80.5,101,-73</points>
<intersection>-80.5 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-73,117,-73</points>
<connection>
<GID>321</GID>
<name>IN_B_3</name></connection>
<intersection>101 0</intersection>
<intersection>117 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-80.5,101,-80.5</points>
<connection>
<GID>297</GID>
<name>OUT_3</name></connection>
<intersection>101 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117,-86.5,117,-73</points>
<intersection>-86.5 4</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>117,-86.5,117.5,-86.5</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>117 3</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-92,100,-72</points>
<intersection>-92 3</intersection>
<intersection>-82.5 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-72,117,-72</points>
<connection>
<GID>321</GID>
<name>IN_B_2</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-82.5,100,-82.5</points>
<connection>
<GID>297</GID>
<name>OUT_2</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>100,-92,117.5,-92</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-97.5,99,-71</points>
<intersection>-97.5 3</intersection>
<intersection>-84.5 2</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-71,117,-71</points>
<connection>
<GID>321</GID>
<name>IN_B_1</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-84.5,99,-84.5</points>
<connection>
<GID>297</GID>
<name>OUT_1</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99,-97.5,117.5,-97.5</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-103,98,-70</points>
<intersection>-103 3</intersection>
<intersection>-86.5 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-70,117,-70</points>
<connection>
<GID>321</GID>
<name>IN_B_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-86.5,98,-86.5</points>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>98,-103,117.5,-103</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-65.5,96.5,-64</points>
<intersection>-65.5 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-64,117,-64</points>
<connection>
<GID>320</GID>
<name>IN_3</name></connection>
<intersection>96.5 0</intersection>
<intersection>116.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-65.5,96.5,-65.5</points>
<connection>
<GID>296</GID>
<name>OUT_3</name></connection>
<intersection>96.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,-106.5,116.5,-64</points>
<intersection>-106.5 4</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>116.5,-106.5,117.5,-106.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>116.5 3</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-0.000100533,235.418,1595,-651.582</PageViewport></page 5>
<page 6>
<PageViewport>0.326052,53.8659,675.516,-321.616</PageViewport>
<gate>
<ID>193</ID>
<type>DD_KEYPAD_HEX</type>
<position>38.5,-28</position>
<output>
<ID>OUT_0</ID>248 </output>
<output>
<ID>OUT_1</ID>247 </output>
<output>
<ID>OUT_2</ID>246 </output>
<output>
<ID>OUT_3</ID>245 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>194</ID>
<type>DD_KEYPAD_HEX</type>
<position>38.5,-43</position>
<output>
<ID>OUT_0</ID>244 </output>
<output>
<ID>OUT_1</ID>243 </output>
<output>
<ID>OUT_2</ID>242 </output>
<output>
<ID>OUT_3</ID>241 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>195</ID>
<type>DD_KEYPAD_HEX</type>
<position>38.5,-57</position>
<output>
<ID>OUT_0</ID>252 </output>
<output>
<ID>OUT_1</ID>251 </output>
<output>
<ID>OUT_2</ID>250 </output>
<output>
<ID>OUT_3</ID>249 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>79,3</position>
<gparam>LABEL_TEXT ALU</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>AA_AND2</type>
<position>77,-46.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_AND2</type>
<position>77,-51.5</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>262 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND2</type>
<position>76.5,-56.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>263 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_AND2</type>
<position>76.5,-61.5</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>264 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND2</type>
<position>76.5,-66.5</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>249 </input>
<output>
<ID>OUT</ID>265 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_AND2</type>
<position>76,-71.5</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_AND2</type>
<position>76,-76.5</position>
<input>
<ID>IN_0</ID>247 </input>
<input>
<ID>IN_1</ID>251 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_AND2</type>
<position>76,-81.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_MUX_2x1</type>
<position>106,-24.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>270 </output>
<input>
<ID>SEL_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_MUX_2x1</type>
<position>105,-31.5</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>267 </input>
<output>
<ID>OUT</ID>271 </output>
<input>
<ID>SEL_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>149,-44.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_MUX_2x1</type>
<position>105.5,-37</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>266 </input>
<output>
<ID>OUT</ID>272 </output>
<input>
<ID>SEL_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>400</ID>
<type>AA_TOGGLE</type>
<position>144,-34</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_MUX_2x1</type>
<position>105.5,-46</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>273 </output>
<input>
<ID>SEL_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>401</ID>
<type>AA_LABEL</type>
<position>157,-33.5</position>
<gparam>LABEL_TEXT Control Signal</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_MUX_2x1</type>
<position>105.5,-52.5</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>264 </input>
<output>
<ID>OUT</ID>274 </output>
<input>
<ID>SEL_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_MUX_2x1</type>
<position>105,-59.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>263 </input>
<output>
<ID>OUT</ID>275 </output>
<input>
<ID>SEL_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_MUX_2x1</type>
<position>105,-66</position>
<input>
<ID>IN_0</ID>254 </input>
<input>
<ID>IN_1</ID>262 </input>
<output>
<ID>OUT</ID>276 </output>
<input>
<ID>SEL_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_MUX_2x1</type>
<position>105,-74.5</position>
<input>
<ID>IN_0</ID>253 </input>
<input>
<ID>IN_1</ID>261 </input>
<output>
<ID>OUT</ID>277 </output>
<input>
<ID>SEL_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_TOGGLE</type>
<position>108.5,-12.5</position>
<output>
<ID>OUT_0</ID>269 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>213</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>137.5,-46</position>
<input>
<ID>IN_0</ID>277 </input>
<input>
<ID>IN_1</ID>276 </input>
<input>
<ID>IN_2</ID>275 </input>
<input>
<ID>IN_3</ID>274 </input>
<input>
<ID>IN_4</ID>273 </input>
<input>
<ID>IN_5</ID>272 </input>
<input>
<ID>IN_6</ID>271 </input>
<input>
<ID>IN_7</ID>270 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 34</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>28,-21</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>29,-49.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>121.5,-12</position>
<gparam>LABEL_TEXT Control Signal</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AE_FULLADDER_4BIT</type>
<position>78,-18.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>247 </input>
<input>
<ID>IN_2</ID>246 </input>
<input>
<ID>IN_3</ID>245 </input>
<input>
<ID>IN_B_0</ID>252 </input>
<input>
<ID>IN_B_1</ID>251 </input>
<input>
<ID>IN_B_2</ID>250 </input>
<input>
<ID>IN_B_3</ID>249 </input>
<output>
<ID>OUT_0</ID>253 </output>
<output>
<ID>OUT_1</ID>254 </output>
<output>
<ID>OUT_2</ID>255 </output>
<output>
<ID>OUT_3</ID>256 </output>
<output>
<ID>carry_out</ID>236 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>191</ID>
<type>AE_FULLADDER_4BIT</type>
<position>77.5,-34.5</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>239 </input>
<input>
<ID>IN_2</ID>238 </input>
<input>
<ID>IN_3</ID>237 </input>
<input>
<ID>IN_B_0</ID>244 </input>
<input>
<ID>IN_B_1</ID>243 </input>
<input>
<ID>IN_B_2</ID>242 </input>
<input>
<ID>IN_B_3</ID>241 </input>
<output>
<ID>OUT_0</ID>257 </output>
<output>
<ID>OUT_1</ID>258 </output>
<output>
<ID>OUT_2</ID>259 </output>
<output>
<ID>OUT_3</ID>260 </output>
<input>
<ID>carry_in</ID>236 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>192</ID>
<type>DD_KEYPAD_HEX</type>
<position>38.5,-14.5</position>
<output>
<ID>OUT_0</ID>240 </output>
<output>
<ID>OUT_1</ID>239 </output>
<output>
<ID>OUT_2</ID>238 </output>
<output>
<ID>OUT_3</ID>237 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>76.5,-26.5,77,-26.5</points>
<connection>
<GID>191</GID>
<name>carry_in</name></connection>
<connection>
<GID>190</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-39.5,58.5,-11.5</points>
<intersection>-39.5 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-39.5,74,-39.5</points>
<connection>
<GID>191</GID>
<name>IN_3</name></connection>
<intersection>58.5 0</intersection>
<intersection>74 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-11.5,58.5,-11.5</points>
<connection>
<GID>192</GID>
<name>OUT_3</name></connection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-45.5,74,-39.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>-39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-38.5,58.5,-13.5</points>
<intersection>-38.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-38.5,74,-38.5</points>
<connection>
<GID>191</GID>
<name>IN_2</name></connection>
<intersection>58.5 0</intersection>
<intersection>74 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-13.5,58.5,-13.5</points>
<connection>
<GID>192</GID>
<name>OUT_2</name></connection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-50.5,74,-38.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>-38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-37.5,58.5,-15.5</points>
<intersection>-37.5 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-37.5,73.5,-37.5</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection>
<intersection>73.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-15.5,58.5,-15.5</points>
<connection>
<GID>192</GID>
<name>OUT_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73.5,-55.5,73.5,-37.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-37.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-36.5,58.5,-17.5</points>
<intersection>-36.5 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-36.5,73.5,-36.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection>
<intersection>73.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-17.5,58.5,-17.5</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73.5,-60.5,73.5,-36.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-40,58.5,-32.5</points>
<intersection>-40 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-32.5,74,-32.5</points>
<connection>
<GID>191</GID>
<name>IN_B_3</name></connection>
<intersection>58.5 0</intersection>
<intersection>74 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-40,58.5,-40</points>
<connection>
<GID>194</GID>
<name>OUT_3</name></connection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-47.5,74,-32.5</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-52.5,58.5,-31.5</points>
<intersection>-52.5 3</intersection>
<intersection>-42 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-31.5,73.5,-31.5</points>
<connection>
<GID>191</GID>
<name>IN_B_2</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-42,58.5,-42</points>
<connection>
<GID>194</GID>
<name>OUT_2</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-52.5,74,-52.5</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-57.5,58.5,-30.5</points>
<intersection>-57.5 3</intersection>
<intersection>-44 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-30.5,73.5,-30.5</points>
<connection>
<GID>191</GID>
<name>IN_B_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-44,58.5,-44</points>
<connection>
<GID>194</GID>
<name>OUT_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-57.5,73.5,-57.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-62.5,58.5,-29.5</points>
<intersection>-62.5 3</intersection>
<intersection>-46 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-29.5,73.5,-29.5</points>
<connection>
<GID>191</GID>
<name>IN_B_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-46,58.5,-46</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-62.5,73.5,-62.5</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-25,58.5,-23.5</points>
<intersection>-25 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-23.5,74,-23.5</points>
<connection>
<GID>190</GID>
<name>IN_3</name></connection>
<intersection>58.5 0</intersection>
<intersection>73.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-25,58.5,-25</points>
<connection>
<GID>193</GID>
<name>OUT_3</name></connection>
<intersection>58.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73.5,-65.5,73.5,-23.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-70.5,58.5,-22.5</points>
<intersection>-70.5 3</intersection>
<intersection>-27 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-22.5,74,-22.5</points>
<connection>
<GID>190</GID>
<name>IN_2</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-27,58.5,-27</points>
<connection>
<GID>193</GID>
<name>OUT_2</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-70.5,73,-70.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-75.5,58.5,-21.5</points>
<intersection>-75.5 3</intersection>
<intersection>-29 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-21.5,74,-21.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-29,58.5,-29</points>
<connection>
<GID>193</GID>
<name>OUT_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-75.5,73,-75.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-80.5,58.5,-20.5</points>
<intersection>-80.5 3</intersection>
<intersection>-31 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-20.5,74,-20.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-31,58.5,-31</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-80.5,73,-80.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-67.5,58.5,-16.5</points>
<intersection>-67.5 3</intersection>
<intersection>-54 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-16.5,74,-16.5</points>
<connection>
<GID>190</GID>
<name>IN_B_3</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-54,58.5,-54</points>
<connection>
<GID>195</GID>
<name>OUT_3</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-67.5,73.5,-67.5</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-72.5,58.5,-15.5</points>
<intersection>-72.5 3</intersection>
<intersection>-56 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-15.5,74,-15.5</points>
<connection>
<GID>190</GID>
<name>IN_B_2</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-56,58.5,-56</points>
<connection>
<GID>195</GID>
<name>OUT_2</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-72.5,73,-72.5</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-77.5,58.5,-14.5</points>
<intersection>-77.5 3</intersection>
<intersection>-58 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-14.5,74,-14.5</points>
<connection>
<GID>190</GID>
<name>IN_B_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-58,58.5,-58</points>
<connection>
<GID>195</GID>
<name>OUT_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-77.5,73,-77.5</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-82.5,58.5,-13.5</points>
<intersection>-82.5 3</intersection>
<intersection>-60 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-13.5,74,-13.5</points>
<connection>
<GID>190</GID>
<name>IN_B_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-60,58.5,-60</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-82.5,73,-82.5</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-75.5,92,-17</points>
<intersection>-75.5 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-75.5,103,-75.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-17,92,-17</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-67,92,-18</points>
<intersection>-67 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-67,103,-67</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-18,92,-18</points>
<connection>
<GID>190</GID>
<name>OUT_1</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-60.5,92.5,-19</points>
<intersection>-60.5 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-60.5,103,-60.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-19,92.5,-19</points>
<connection>
<GID>190</GID>
<name>OUT_2</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-53.5,92.5,-20</points>
<intersection>-53.5 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-53.5,103.5,-53.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-20,92.5,-20</points>
<connection>
<GID>190</GID>
<name>OUT_3</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-47,92.5,-33</points>
<intersection>-47 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-47,103.5,-47</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-33,92.5,-33</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-38,92.5,-34</points>
<intersection>-38 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-38,103.5,-38</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-34,92.5,-34</points>
<connection>
<GID>191</GID>
<name>OUT_1</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-35,92.5,-32.5</points>
<intersection>-35 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-32.5,103,-32.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-35,92.5,-35</points>
<connection>
<GID>191</GID>
<name>OUT_2</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-36,92.5,-25.5</points>
<intersection>-36 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-25.5,104,-25.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-36,92.5,-36</points>
<connection>
<GID>191</GID>
<name>OUT_3</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-73.5,91.5,-46.5</points>
<intersection>-73.5 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-73.5,103,-73.5</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80,-46.5,91.5,-46.5</points>
<connection>
<GID>196</GID>
<name>OUT</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-65,91.5,-51.5</points>
<intersection>-65 1</intersection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-65,103,-65</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80,-51.5,91.5,-51.5</points>
<connection>
<GID>197</GID>
<name>OUT</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-58.5,91,-56.5</points>
<intersection>-58.5 1</intersection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91,-58.5,103,-58.5</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>91 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79.5,-56.5,91,-56.5</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-61.5,91.5,-51.5</points>
<intersection>-61.5 2</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-51.5,103.5,-51.5</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79.5,-61.5,91.5,-61.5</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-66.5,91.5,-45</points>
<intersection>-66.5 2</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-45,103.5,-45</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79.5,-66.5,91.5,-66.5</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-71.5,91,-36</points>
<intersection>-71.5 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91,-36,103.5,-36</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>91 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,-71.5,91,-71.5</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-76.5,91.5,-30.5</points>
<intersection>-76.5 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-30.5,103,-30.5</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,-76.5,91.5,-76.5</points>
<connection>
<GID>202</GID>
<name>OUT</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-81.5,91.5,-23.5</points>
<intersection>-81.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-23.5,104,-23.5</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,-81.5,91.5,-81.5</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-34.5,105,-12.5</points>
<connection>
<GID>205</GID>
<name>SEL_0</name></connection>
<intersection>-34.5 3</intersection>
<intersection>-22 9</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-12.5,106.5,-12.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105,-34.5,105.5,-34.5</points>
<connection>
<GID>206</GID>
<name>SEL_0</name></connection>
<intersection>105 0</intersection>
<intersection>105.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>105.5,-57,105.5,-34.5</points>
<connection>
<GID>207</GID>
<name>SEL_0</name></connection>
<connection>
<GID>208</GID>
<name>SEL_0</name></connection>
<intersection>-57 6</intersection>
<intersection>-34.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>105,-57,105.5,-57</points>
<connection>
<GID>209</GID>
<name>SEL_0</name></connection>
<intersection>105 7</intersection>
<intersection>105.5 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>105,-72,105,-57</points>
<connection>
<GID>210</GID>
<name>SEL_0</name></connection>
<connection>
<GID>211</GID>
<name>SEL_0</name></connection>
<intersection>-57 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>105,-22,106,-22</points>
<connection>
<GID>204</GID>
<name>SEL_0</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-42,130.5,-24.5</points>
<intersection>-42 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-42,132.5,-42</points>
<connection>
<GID>213</GID>
<name>IN_7</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108,-24.5,130.5,-24.5</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-43,129,-31.5</points>
<intersection>-43 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129,-43,132.5,-43</points>
<connection>
<GID>213</GID>
<name>IN_6</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107,-31.5,129,-31.5</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-44,120,-37</points>
<intersection>-44 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-44,132.5,-44</points>
<connection>
<GID>213</GID>
<name>IN_5</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-37,120,-37</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-46,120,-45</points>
<intersection>-46 2</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-45,132.5,-45</points>
<connection>
<GID>213</GID>
<name>IN_4</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-46,120,-46</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-52.5,120,-46</points>
<intersection>-52.5 2</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-46,132.5,-46</points>
<connection>
<GID>213</GID>
<name>IN_3</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-52.5,120,-52.5</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-59.5,119.5,-47</points>
<intersection>-59.5 2</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-47,132.5,-47</points>
<connection>
<GID>213</GID>
<name>IN_2</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107,-59.5,119.5,-59.5</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-66,119.5,-48</points>
<intersection>-66 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-48,132.5,-48</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107,-66,119.5,-66</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-74.5,119.5,-49</points>
<intersection>-74.5 2</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-49,132.5,-49</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107,-74.5,119.5,-74.5</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>-0.000100533,235.418,1595,-651.582</PageViewport></page 7>
<page 8>
<PageViewport>-0.000100533,235.418,1595,-651.582</PageViewport></page 8>
<page 9>
<PageViewport>-0.000100533,235.418,1595,-651.582</PageViewport></page 9></circuit>